magic
tech sky130A
magscale 1 2
timestamp 1634488599
<< error_s >>
rect 298 981 333 1015
rect 299 962 333 981
rect 129 913 187 919
rect 129 879 141 913
rect 129 873 187 879
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 318 583 333 962
rect 352 928 387 962
rect 667 928 702 962
rect 352 583 386 928
rect 668 909 702 928
rect 498 860 556 866
rect 498 826 510 860
rect 498 820 556 826
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 352 549 367 583
rect 687 530 702 909
rect 721 875 756 909
rect 1036 875 1071 909
rect 721 530 755 875
rect 1037 856 1071 875
rect 867 807 925 813
rect 867 773 879 807
rect 867 767 925 773
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 721 496 736 530
rect 1056 477 1071 856
rect 1090 822 1125 856
rect 1405 822 1440 856
rect 1090 477 1124 822
rect 1406 803 1440 822
rect 1236 754 1294 760
rect 1236 720 1248 754
rect 1236 714 1294 720
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1425 424 1440 803
rect 1459 769 1494 803
rect 1774 769 1809 803
rect 1459 424 1493 769
rect 1775 750 1809 769
rect 1605 701 1663 707
rect 1605 667 1617 701
rect 1605 661 1663 667
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1794 371 1809 750
rect 1828 716 1863 750
rect 2143 716 2178 750
rect 1828 371 1862 716
rect 2144 697 2178 716
rect 2530 697 2583 698
rect 1974 648 2032 654
rect 1974 614 1986 648
rect 1974 608 2032 614
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1828 337 1843 371
rect 2163 318 2178 697
rect 2197 663 2232 697
rect 2512 663 2583 697
rect 2197 318 2231 663
rect 2513 662 2583 663
rect 2530 628 2601 662
rect 2921 628 2956 662
rect 2343 595 2401 601
rect 2343 561 2355 595
rect 2343 555 2401 561
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2530 265 2600 628
rect 2922 609 2956 628
rect 2730 560 2792 566
rect 2730 526 2742 560
rect 2730 520 2792 526
rect 2730 348 2792 354
rect 2730 314 2742 348
rect 2730 308 2792 314
rect 2530 229 2583 265
rect 2941 212 2956 609
rect 2975 575 3010 609
rect 3330 575 3365 609
rect 2975 212 3009 575
rect 3331 556 3365 575
rect 3139 507 3201 513
rect 3139 473 3151 507
rect 3139 467 3201 473
rect 3139 295 3201 301
rect 3139 261 3151 295
rect 3139 255 3201 261
rect 2975 178 2990 212
rect 3350 159 3365 556
rect 3384 522 3419 556
rect 3739 522 3774 556
rect 3384 159 3418 522
rect 3740 503 3774 522
rect 3548 454 3610 460
rect 3548 420 3560 454
rect 3548 414 3610 420
rect 3548 242 3610 248
rect 3548 208 3560 242
rect 3548 202 3610 208
rect 3384 125 3399 159
rect 3759 106 3774 503
rect 3793 469 3828 503
rect 4148 469 4183 503
rect 3793 106 3827 469
rect 4149 450 4183 469
rect 3957 401 4019 407
rect 3957 367 3969 401
rect 3957 361 4019 367
rect 3957 189 4019 195
rect 3957 155 3969 189
rect 3957 149 4019 155
rect 3793 72 3808 106
rect 4168 53 4183 450
rect 4202 416 4237 450
rect 4557 416 4592 450
rect 4202 53 4236 416
rect 4558 397 4592 416
rect 4366 348 4428 354
rect 4366 314 4378 348
rect 4366 308 4428 314
rect 4366 136 4428 142
rect 4366 102 4378 136
rect 4366 96 4428 102
rect 4202 19 4217 53
rect 4577 0 4592 397
rect 4611 363 4646 397
rect 4966 363 5001 380
rect 4611 0 4645 363
rect 4967 362 5001 363
rect 4967 326 5037 362
rect 4775 295 4837 301
rect 4775 261 4787 295
rect 4984 292 5055 326
rect 5335 292 5370 326
rect 4775 255 4837 261
rect 4775 83 4837 89
rect 4775 49 4787 83
rect 4775 43 4837 49
rect 4611 -34 4626 0
rect 4984 -53 5054 292
rect 5336 273 5370 292
rect 5722 273 5775 274
rect 5166 224 5224 230
rect 5166 190 5178 224
rect 5166 184 5224 190
rect 5166 30 5224 36
rect 5166 -4 5178 30
rect 5166 -10 5224 -4
rect 4984 -89 5037 -53
rect 5355 -106 5370 273
rect 5389 239 5424 273
rect 5704 239 5775 273
rect 5389 -106 5423 239
rect 5705 238 5775 239
rect 5722 204 5793 238
rect 6113 204 6148 221
rect 5535 171 5593 177
rect 5535 137 5547 171
rect 5535 131 5593 137
rect 5535 -23 5593 -17
rect 5535 -57 5547 -23
rect 5535 -63 5593 -57
rect 5389 -140 5404 -106
rect 5722 -159 5792 204
rect 6114 203 6148 204
rect 6114 167 6184 203
rect 5922 136 5984 142
rect 5922 102 5934 136
rect 6131 133 6202 167
rect 6482 133 6517 167
rect 5922 96 5984 102
rect 5922 -76 5984 -70
rect 5922 -110 5934 -76
rect 5922 -116 5984 -110
rect 5722 -195 5775 -159
rect 6131 -212 6201 133
rect 6483 114 6517 133
rect 6313 65 6371 71
rect 6313 31 6325 65
rect 6313 25 6371 31
rect 6313 -129 6371 -123
rect 6313 -163 6325 -129
rect 6313 -169 6371 -163
rect 6131 -248 6184 -212
rect 6502 -265 6517 114
rect 6536 80 6571 114
rect 6536 -265 6570 80
rect 6682 12 6740 18
rect 6682 -22 6694 12
rect 6682 -28 6740 -22
rect 6682 -182 6740 -176
rect 6682 -216 6694 -182
rect 6682 -222 6740 -216
rect 6536 -299 6551 -265
rect 6922 -318 6940 168
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  X1
timestamp 1634488599
transform 1 0 158 0 1 799
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  X2
timestamp 1634488599
transform 1 0 527 0 1 746
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  X3
timestamp 1634488599
transform 1 0 896 0 1 693
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  X4
timestamp 1634488599
transform 1 0 1265 0 1 640
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  X5
timestamp 1634488599
transform 1 0 1634 0 1 587
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  X6
timestamp 1634488599
transform 1 0 2003 0 1 534
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  X7
timestamp 1634488599
transform 1 0 2372 0 1 481
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_lvt_EM43P7  X8
timestamp 1634488599
transform 1 0 2761 0 1 437
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_EM43P7  X9
timestamp 1634488599
transform 1 0 3170 0 1 384
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_EM43P7  X10
timestamp 1634488599
transform 1 0 3579 0 1 331
box -231 -261 231 261
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ0
timestamp 1634257435
transform 1 0 6896 0 1 -380
box 26 26 770 795
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  Xf
timestamp 1634488599
transform 1 0 6711 0 1 -102
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  Xe
timestamp 1634488599
transform 1 0 6342 0 1 -49
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_lvt_EM43P7  Xd
timestamp 1634488599
transform 1 0 5953 0 1 13
box -231 -261 231 261
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  Xc
timestamp 1634488599
transform 1 0 5564 0 1 57
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_L7T3GD  Xb
timestamp 1634488599
transform 1 0 5195 0 1 110
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_lvt_EM43P7  Xa
timestamp 1634488599
transform 1 0 4806 0 1 172
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_EM43P7  X12
timestamp 1634488599
transform 1 0 4397 0 1 225
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_EM43P7  X11
timestamp 1634488599
transform 1 0 3988 0 1 278
box -231 -261 231 261
<< end >>
