magic
tech sky130A
magscale 1 2
timestamp 1634541323
<< nmoslvt >>
rect -229 -800 -29 800
rect 29 -800 229 800
<< ndiff >>
rect -287 788 -229 800
rect -287 -788 -275 788
rect -241 -788 -229 788
rect -287 -800 -229 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 229 788 287 800
rect 229 -788 241 788
rect 275 -788 287 788
rect 229 -800 287 -788
<< ndiffc >>
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
<< poly >>
rect -187 872 -71 888
rect -187 855 -171 872
rect -229 838 -171 855
rect -87 855 -71 872
rect 71 872 187 888
rect 71 855 87 872
rect -87 838 -29 855
rect -229 800 -29 838
rect 29 838 87 855
rect 171 855 187 872
rect 171 838 229 855
rect 29 800 229 838
rect -229 -838 -29 -800
rect -229 -855 -171 -838
rect -187 -872 -171 -855
rect -87 -855 -29 -838
rect 29 -838 229 -800
rect 29 -855 87 -838
rect -87 -872 -71 -855
rect -187 -888 -71 -872
rect 71 -872 87 -855
rect 171 -855 229 -838
rect 171 -872 187 -855
rect 71 -888 187 -872
<< polycont >>
rect -171 838 -87 872
rect 87 838 171 872
rect -171 -872 -87 -838
rect 87 -872 171 -838
<< locali >>
rect -187 838 -171 872
rect -87 838 -71 872
rect 71 838 87 872
rect 171 838 187 872
rect -275 788 -241 804
rect -275 -804 -241 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 241 788 275 804
rect 241 -804 275 -788
rect -187 -872 -171 -838
rect -87 -872 -71 -838
rect 71 -872 87 -838
rect 171 -872 187 -838
<< viali >>
rect -171 838 -87 872
rect 87 838 171 872
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect -171 -872 -87 -838
rect 87 -872 171 -838
<< metal1 >>
rect -183 872 -75 878
rect -183 838 -171 872
rect -87 838 -75 872
rect -183 832 -75 838
rect 75 872 183 878
rect 75 838 87 872
rect 171 838 183 872
rect 75 832 183 838
rect -281 788 -235 800
rect -281 -788 -275 788
rect -241 -788 -235 788
rect -281 -800 -235 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 235 788 281 800
rect 235 -788 241 788
rect 275 -788 281 788
rect 235 -800 281 -788
rect -183 -838 -75 -832
rect -183 -872 -171 -838
rect -87 -872 -75 -838
rect -183 -878 -75 -872
rect 75 -838 183 -832
rect 75 -872 87 -838
rect 171 -872 183 -838
rect 75 -878 183 -872
<< labels >>
flabel metal1 -23 -800 -17 800 0 FreeSans 160 0 0 0 S$
flabel metal1 17 -800 23 800 0 FreeSans 160 0 0 0 S$
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 8 l 1 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
