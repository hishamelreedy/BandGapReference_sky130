magic
tech sky130A
magscale 1 2
timestamp 1634815686
<< nwell >>
rect 1790 4006 2036 4040
rect 1790 4002 2048 4006
rect 1790 1334 2036 4002
rect 5532 3578 5612 3758
rect 5492 3502 5636 3578
rect 5520 1504 5612 3502
rect 6072 3358 6550 3952
rect 5488 1402 5638 1504
rect 5880 1428 6624 3358
rect 2030 1146 2048 1296
rect 5532 1118 5612 1402
rect 2846 256 2950 388
<< nsubdiff >>
rect 1844 3530 1988 3578
rect 1844 3502 1872 3530
rect 1840 1454 1872 1504
rect 1952 3502 1988 3530
rect 5492 3530 5636 3578
rect 5492 3502 5520 3530
rect 1952 1454 1990 1504
rect 1840 1402 1990 1454
rect 5488 1454 5520 1504
rect 5600 3502 5636 3530
rect 5600 1454 5638 1504
rect 5488 1402 5638 1454
<< nsubdiffcont >>
rect 1872 1454 1952 3530
rect 5520 1454 5600 3530
<< locali >>
rect 1814 3674 2010 3710
rect 1814 3586 1842 3674
rect 1988 3586 2010 3674
rect 1814 3576 2010 3586
rect 5462 3674 5658 3710
rect 5462 3586 5490 3674
rect 5636 3586 5658 3674
rect 5462 3576 5658 3586
rect 1838 3540 1990 3576
rect 5486 3540 5638 3576
rect 1844 3530 1988 3540
rect 1844 3502 1872 3530
rect 1840 1454 1872 1504
rect 1952 3502 1988 3530
rect 5492 3530 5636 3540
rect 5492 3502 5520 3530
rect 1952 1454 1990 1504
rect 1840 1402 1990 1454
rect 5488 1454 5520 1504
rect 5600 3502 5636 3530
rect 5600 1454 5638 1504
rect 5488 1402 5638 1454
<< viali >>
rect 1842 3586 1988 3674
rect 5490 3586 5636 3674
<< metal1 >>
rect 1848 3964 1974 3976
rect 1848 3898 1866 3964
rect 1952 3898 1974 3964
rect -4826 3858 -4470 3876
rect -4826 3808 -4758 3858
rect -4830 3732 -4758 3808
rect -4826 3658 -4758 3732
rect -4568 3808 -4470 3858
rect -4568 3732 -518 3808
rect -4568 3658 -4470 3732
rect 1848 3710 1974 3898
rect 5496 3964 5622 3976
rect 5496 3898 5514 3964
rect 5600 3898 5622 3964
rect 5496 3710 5622 3898
rect -4826 3602 -4470 3658
rect 1814 3674 2010 3710
rect 1814 3586 1842 3674
rect 1988 3586 2010 3674
rect 1814 3576 2010 3586
rect 5462 3674 5658 3710
rect 5462 3586 5490 3674
rect 5636 3586 5658 3674
rect 5462 3576 5658 3586
rect -4792 3110 -4436 3146
rect -4792 2910 -4726 3110
rect -4536 3042 -4436 3110
rect -4536 2966 -436 3042
rect -4536 2910 -4436 2966
rect -4792 2872 -4436 2910
rect -4810 1480 -4414 1534
rect -4810 1174 -4748 1480
rect -4488 1174 -4414 1480
rect -4810 1154 -4414 1174
rect -1294 932 -1076 956
rect 1656 946 1878 960
rect 1656 764 3018 946
rect 1656 516 1878 764
rect -2682 422 1878 516
rect 1656 346 1878 422
rect -4664 -562 -4418 -522
rect -4664 -762 -4636 -562
rect -4446 -634 -4418 -562
rect -4446 -664 -528 -634
rect -4446 -762 -4418 -664
rect -4664 -796 -4418 -762
rect -4680 -1250 -4434 -1214
rect -4680 -1362 -4648 -1250
rect -4684 -1392 -4648 -1362
rect -4680 -1450 -4648 -1392
rect -4458 -1362 -4434 -1250
rect -4458 -1392 -760 -1362
rect -4458 -1450 -4434 -1392
rect -4680 -1488 -4434 -1450
rect -4714 -1970 -4468 -1952
rect -4714 -2170 -4692 -1970
rect -4502 -2096 -4468 -1970
rect -4502 -2126 -782 -2096
rect -4502 -2170 -4468 -2126
rect -4714 -2226 -4468 -2170
rect -4708 -2728 -4462 -2700
rect -4708 -2928 -4676 -2728
rect -4486 -2852 -4462 -2728
rect -4486 -2882 -666 -2852
rect -4486 -2928 -4462 -2882
rect -4708 -2974 -4462 -2928
rect 7932 -3096 8292 -3046
rect 7932 -3168 7964 -3096
rect 1268 -3220 7964 -3168
rect 7932 -3288 7964 -3220
rect 8240 -3288 8292 -3096
rect 7932 -3344 8292 -3288
rect -4212 -5932 -3457 -5872
rect -4640 -6458 -4408 -6456
rect -4644 -6474 -4408 -6458
rect -4644 -6564 -4578 -6474
rect -4444 -6508 -4408 -6474
rect -4444 -6510 -544 -6508
rect -4444 -6540 -484 -6510
rect -4444 -6564 -4408 -6540
rect -4644 -6582 -4408 -6564
rect -4644 -6584 -4412 -6582
rect -4628 -7202 -4396 -7190
rect -4628 -7292 -4556 -7202
rect -4422 -7260 -4396 -7202
rect -4422 -7290 -494 -7260
rect -4422 -7292 -4396 -7290
rect -4628 -7316 -4396 -7292
<< via1 >>
rect 1866 3898 1952 3964
rect -4758 3658 -4568 3858
rect 5514 3898 5600 3964
rect -4726 2910 -4536 3110
rect -4748 1174 -4488 1480
rect -4636 -762 -4446 -562
rect -4648 -1450 -4458 -1250
rect -4692 -2170 -4502 -1970
rect -4676 -2928 -4486 -2728
rect 7964 -3288 8240 -3096
rect -4578 -6564 -4444 -6474
rect -4556 -7292 -4422 -7202
<< metal2 >>
rect -5144 4972 8554 5464
rect -5240 3858 -4410 4070
rect 1790 3964 2015 4026
rect 1790 3898 1866 3964
rect 1952 3898 2015 3964
rect 1790 3884 2015 3898
rect 2428 3860 2692 4972
rect 3494 3886 3758 4972
rect 4322 3886 4586 4972
rect 5024 3886 5288 4972
rect -5240 3658 -4758 3858
rect -4568 3658 -4410 3858
rect -5240 3110 -4410 3658
rect -5240 2910 -4726 3110
rect -4536 2910 -4410 3110
rect -5240 1480 -4410 2910
rect -5240 1174 -4748 1480
rect -4488 1174 -4410 1480
rect -5240 -562 -4410 1174
rect 4758 412 6192 418
rect 2836 240 2952 396
rect 3000 344 3108 394
rect 3000 258 3022 344
rect 3090 258 3108 344
rect 2868 -108 2932 240
rect 3000 226 3108 258
rect 3776 206 3892 234
rect 3776 120 3798 206
rect 3866 120 3892 206
rect 3776 78 3892 120
rect 3998 180 4092 242
rect 4758 230 6198 412
rect 3998 174 4684 180
rect 3998 76 4804 174
rect 2868 -184 3466 -108
rect -5240 -762 -4636 -562
rect -4446 -762 -4410 -562
rect 3286 -634 3460 -184
rect 4548 -754 4804 76
rect -5240 -1250 -4410 -762
rect 5902 -844 6198 230
rect -5240 -1450 -4648 -1250
rect -4458 -1450 -4410 -1250
rect -5240 -1970 -4410 -1450
rect 6836 -1548 8550 -1214
rect -5240 -2170 -4692 -1970
rect -4502 -2170 -4410 -1970
rect -5240 -2728 -4410 -2170
rect -5240 -2928 -4676 -2728
rect -4486 -2928 -4410 -2728
rect -5240 -6474 -4410 -2928
rect 7936 -3096 8408 -2632
rect 7936 -3288 7964 -3096
rect 8240 -3288 8408 -3096
rect -5240 -6564 -4578 -6474
rect -4444 -6564 -4410 -6474
rect -5240 -7202 -4410 -6564
rect -5240 -7292 -4556 -7202
rect -4422 -7292 -4410 -7202
rect -5240 -8274 -4410 -7292
rect -274 -8274 -136 -6058
rect 7936 -8274 8408 -3288
rect -5240 -8332 8460 -8274
rect -5238 -8766 8460 -8332
<< via2 >>
rect 3442 970 3510 1056
rect 3022 258 3090 344
rect 3798 120 3866 206
rect 2020 -932 2088 -846
rect 6936 -984 7004 -898
rect 592 -1474 660 -1388
<< metal3 >>
rect 3428 1056 7090 1074
rect 3428 970 3442 1056
rect 3510 970 7090 1056
rect 3428 940 7090 970
rect 3002 344 3106 358
rect 3002 258 3022 344
rect 3090 258 3106 344
rect 3002 234 3106 258
rect 3014 176 3088 234
rect 3786 206 3880 224
rect 3014 172 3086 176
rect 1992 -268 2900 -264
rect 3016 -268 3086 172
rect 3786 120 3798 206
rect 3866 120 3880 206
rect 3786 112 3880 120
rect 3786 92 3882 112
rect 3790 6 3882 92
rect 1992 -328 3086 -268
rect 1992 -332 3084 -328
rect 1992 -846 2118 -332
rect 1992 -932 2020 -846
rect 2088 -932 2118 -846
rect 1992 -978 2118 -932
rect 3792 -1316 3882 6
rect 6898 -898 7090 940
rect 6898 -984 6936 -898
rect 7004 -984 7090 -898
rect 6898 -1028 7090 -984
rect 530 -1388 3884 -1316
rect 530 -1474 592 -1388
rect 660 -1474 3884 -1388
rect 530 -1538 3884 -1474
use pmos_mirror  pmos_mirror_0
timestamp 1634671827
transform 1 0 4180 0 1 2174
box -4180 -2174 3034 2473
use PDN  PDN_0
timestamp 1634813859
transform 1 0 6158 0 1 -4980
box -11370 -3742 1046 9021
<< labels >>
flabel metal2 6836 -1548 8550 -1214 0 FreeSans 1600 0 0 0 VBGP
flabel metal2 -5144 4972 8554 5464 0 FreeSans 1600 0 0 0 VDD
flabel metal2 -5238 -8766 8460 -8274 0 FreeSans 1600 0 0 0 AGND
<< end >>
