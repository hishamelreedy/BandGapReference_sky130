magic
tech sky130A
timestamp 1635333008
<< psubdiff >>
rect -447 7471 -107 7475
rect -447 7453 51 7471
rect 7009 7470 7329 7483
rect 6876 7467 7329 7470
rect 6873 7453 7329 7467
rect -447 7166 36 7453
rect 6888 7166 7329 7453
rect -447 7135 51 7166
rect 6873 7157 7329 7166
rect 6876 7151 7329 7157
rect 7009 7139 7329 7151
rect -447 7075 -107 7135
rect -447 7040 -424 7075
rect -444 223 -424 314
rect -137 7040 -107 7075
rect 7009 7066 7041 7139
rect -137 223 -118 314
rect -444 -19 -118 223
rect 7026 287 7041 324
rect 7328 7066 7329 7139
rect 7328 287 7346 324
rect -458 -44 30 -19
rect 7026 -23 7346 287
rect 6795 -44 7346 -23
rect -458 -331 -8 -44
rect 6844 -331 7346 -44
rect -458 -367 30 -331
rect 6795 -349 7346 -331
rect 7026 -360 7346 -349
<< psubdiffcont >>
rect 36 7166 6888 7453
rect -424 223 -137 7075
rect 7041 287 7328 7139
rect -8 -331 6844 -44
<< locali >>
rect -447 7471 -107 7475
rect -447 7453 51 7471
rect 6871 7470 6897 7471
rect 7009 7470 7329 7483
rect 6871 7453 7329 7470
rect -447 7166 36 7453
rect 6888 7166 7329 7453
rect -447 7135 51 7166
rect 6871 7151 7329 7166
rect 6871 7150 6897 7151
rect 7009 7139 7329 7151
rect -447 7075 -107 7135
rect -447 7040 -424 7075
rect -444 223 -424 314
rect -137 7040 -107 7075
rect 7009 7066 7041 7139
rect 7328 7066 7329 7139
rect -137 223 -118 314
rect -444 -19 -118 223
rect 7026 287 7041 324
rect 7328 287 7346 324
rect -458 -44 30 -19
rect 7026 -23 7346 287
rect 6795 -44 7346 -23
rect -458 -331 -8 -44
rect 6844 -331 7346 -44
rect -458 -367 30 -331
rect 6795 -349 7346 -331
rect 7026 -360 7346 -349
<< viali >>
rect 280 7248 376 7349
rect 539 7248 635 7349
rect 801 7248 897 7349
rect 1048 7251 1144 7352
rect 4400 7261 4496 7362
rect 4743 7261 4839 7362
rect 5098 7273 5194 7374
rect 7136 6128 7232 6229
rect 7128 5851 7224 5952
rect 7120 5542 7216 5643
rect 7076 2240 7295 2436
rect 7072 1865 7291 2061
rect 214 -286 433 -90
<< metal1 >>
rect 100 7353 2208 7542
rect 100 7352 1300 7353
rect 100 7349 1048 7352
rect 100 7248 280 7349
rect 376 7248 539 7349
rect 635 7248 801 7349
rect 897 7251 1048 7349
rect 1144 7252 1300 7352
rect 1396 7352 2208 7353
rect 1396 7252 1552 7352
rect 1144 7251 1552 7252
rect 1648 7251 1801 7352
rect 1897 7251 2208 7352
rect 897 7248 2208 7251
rect 100 7143 2208 7248
rect 4254 7374 6672 7524
rect 4254 7362 5098 7374
rect 4254 7261 4400 7362
rect 4496 7261 4743 7362
rect 4839 7273 5098 7362
rect 5194 7273 6672 7374
rect 4839 7261 6672 7273
rect 4254 7126 6672 7261
rect -1348 339 -145 6344
rect 6930 6229 7397 6390
rect 6930 6128 7136 6229
rect 7232 6128 7397 6229
rect 6930 5952 7397 6128
rect 6930 5851 7128 5952
rect 7224 5851 7397 5952
rect 6930 5643 7397 5851
rect 6930 5542 7120 5643
rect 7216 5542 7397 5643
rect 6930 4655 7397 5542
rect 6932 2436 7409 2549
rect 6932 2240 7076 2436
rect 7295 2240 7409 2436
rect 6932 2061 7409 2240
rect 6932 1865 7072 2061
rect 7291 1865 7409 2061
rect 6932 689 7409 1865
rect 33 -90 6840 158
rect 33 -286 214 -90
rect 433 -286 6840 -90
rect 33 -1075 6840 -286
<< via1 >>
rect 280 7248 376 7349
rect 539 7248 635 7349
rect 801 7248 897 7349
rect 1048 7251 1144 7352
rect 1300 7252 1396 7353
rect 1552 7251 1648 7352
rect 1801 7251 1897 7352
rect 4400 7261 4496 7362
rect 4743 7261 4839 7362
rect 5098 7273 5194 7374
rect 7136 6128 7232 6229
rect 7128 5851 7224 5952
rect 7120 5542 7216 5643
rect 7076 2240 7295 2436
rect 7072 1865 7291 2061
rect 214 -286 433 -90
<< metal2 >>
rect 2982 8013 3860 8055
rect 2982 7673 3152 8013
rect 3620 7673 3860 8013
rect 105 7353 2156 7420
rect 105 7352 1300 7353
rect 105 7349 1048 7352
rect 105 7248 280 7349
rect 376 7248 539 7349
rect 635 7248 801 7349
rect 897 7251 1048 7349
rect 1144 7252 1300 7352
rect 1396 7352 2156 7353
rect 1396 7252 1552 7352
rect 1144 7251 1552 7252
rect 1648 7251 1801 7352
rect 1897 7251 2156 7352
rect 897 7248 2156 7251
rect 105 7203 2156 7248
rect 2982 7036 3860 7673
rect 4277 7374 6563 7446
rect 4277 7362 5098 7374
rect 4277 7261 4400 7362
rect 4496 7261 4743 7362
rect 4839 7273 5098 7362
rect 5194 7273 6563 7374
rect 4839 7261 6563 7273
rect 4277 7227 6563 7261
rect -1348 339 -145 6344
rect 6993 6229 7350 6358
rect 6993 6128 7136 6229
rect 7232 6128 7350 6229
rect 6993 5952 7350 6128
rect 6993 5851 7128 5952
rect 7224 5851 7350 5952
rect 6993 5643 7350 5851
rect 6993 5542 7120 5643
rect 7216 5542 7350 5643
rect 6993 4702 7350 5542
rect 6041 3903 7835 4104
rect 6023 3819 7835 3903
rect 6023 3548 7497 3819
rect 7735 3548 7835 3819
rect 6023 3456 7835 3548
rect 6041 3230 7835 3456
rect 7016 2436 7351 2496
rect 7016 2240 7076 2436
rect 7295 2240 7351 2436
rect 7016 2061 7351 2240
rect 7016 1865 7072 2061
rect 7291 1865 7351 2061
rect 7016 713 7351 1865
rect 33 -90 6840 158
rect 33 -286 214 -90
rect 433 -286 6840 -90
rect 33 -1075 6840 -286
<< via2 >>
rect 3152 7673 3620 8013
rect 280 7248 376 7349
rect 539 7248 635 7349
rect 801 7248 897 7349
rect 1048 7251 1144 7352
rect 1300 7252 1396 7353
rect 1552 7251 1648 7352
rect 1801 7251 1897 7352
rect 4400 7261 4496 7362
rect 4743 7261 4839 7362
rect 5098 7273 5194 7374
rect 7136 6128 7232 6229
rect 7128 5851 7224 5952
rect 7120 5542 7216 5643
rect 7497 3548 7735 3819
rect 7076 2240 7295 2436
rect 7072 1865 7291 2061
rect 214 -286 433 -90
<< metal3 >>
rect 2968 8013 3860 8679
rect 2968 7673 3152 8013
rect 3620 7673 3860 8013
rect 2968 7616 3860 7673
rect 95 7353 2183 7589
rect 95 7352 1300 7353
rect 95 7349 1048 7352
rect 95 7248 280 7349
rect 376 7248 539 7349
rect 635 7248 801 7349
rect 897 7251 1048 7349
rect 1144 7252 1300 7352
rect 1396 7352 2183 7353
rect 1396 7252 1552 7352
rect 1144 7251 1552 7252
rect 1648 7251 1801 7352
rect 1897 7251 2183 7352
rect 897 7248 2183 7251
rect 95 7189 2183 7248
rect 4262 7401 6579 7742
rect 4262 7386 6088 7401
rect 4262 7378 5613 7386
rect 4262 7374 5398 7378
rect 4262 7362 5098 7374
rect 4262 7261 4400 7362
rect 4496 7261 4743 7362
rect 4839 7273 5098 7362
rect 5194 7277 5398 7374
rect 5494 7285 5613 7378
rect 5709 7362 6088 7386
rect 5709 7285 5890 7362
rect 5494 7277 5890 7285
rect 5194 7273 5890 7277
rect 4839 7261 5890 7273
rect 5986 7300 6088 7362
rect 6184 7389 6579 7401
rect 6184 7300 6272 7389
rect 5986 7288 6272 7300
rect 6368 7288 6579 7389
rect 5986 7261 6579 7288
rect 4262 7227 6579 7261
rect -1348 5998 -145 6344
rect -1348 5897 -327 5998
rect -231 5897 -145 5998
rect -1348 5205 -145 5897
rect -1348 5104 -327 5205
rect -231 5104 -145 5205
rect -1348 4395 -145 5104
rect 7080 6229 8221 6319
rect 7080 6128 7136 6229
rect 7232 6128 8221 6229
rect 7080 5952 8221 6128
rect 7080 5851 7128 5952
rect 7224 5851 8221 5952
rect 7080 5643 8221 5851
rect 7080 5542 7120 5643
rect 7216 5542 8221 5643
rect 7080 5358 8221 5542
rect 7080 5257 7120 5358
rect 7216 5257 8221 5358
rect 7080 5120 8221 5257
rect 7080 5019 7104 5120
rect 7200 5019 8221 5120
rect 7080 4994 8221 5019
rect 7080 4893 7120 4994
rect 7216 4893 8221 4994
rect 7080 4718 8221 4893
rect -1348 4294 -343 4395
rect -247 4294 -145 4395
rect -1348 3750 -145 4294
rect -1348 3649 -310 3750
rect -214 3649 -145 3750
rect -1348 3287 -145 3649
rect -1348 3186 -310 3287
rect -214 3186 -145 3287
rect 7489 3819 8208 4085
rect 7489 3548 7497 3819
rect 7735 3548 8208 3819
rect 7489 3240 8208 3548
rect -1348 2775 -145 3186
rect -1348 2674 -294 2775
rect -198 2674 -145 2775
rect -1348 2262 -145 2674
rect -1348 2161 -310 2262
rect -214 2161 -145 2262
rect -1348 1783 -145 2161
rect -1348 1682 -310 1783
rect -214 1682 -145 1783
rect -1348 1303 -145 1682
rect -1348 1202 -277 1303
rect -181 1202 -145 1303
rect -1348 791 -145 1202
rect -1348 690 -310 791
rect -214 690 -145 791
rect 7048 2436 7503 2448
rect 7048 2240 7076 2436
rect 7295 2240 7503 2436
rect 7048 2061 7503 2240
rect 7048 1865 7072 2061
rect 7291 1865 7503 2061
rect 7048 1693 7503 1865
rect 7048 1497 7080 1693
rect 7299 1497 7503 1693
rect 7048 1417 7503 1497
rect 7048 1221 7084 1417
rect 7303 1221 7503 1417
rect 7048 1173 7503 1221
rect 7048 977 7092 1173
rect 7311 977 7503 1173
rect 7048 737 7503 977
rect -1348 339 -145 690
rect 33 -8 6840 158
rect 33 -24 4933 -8
rect 33 -40 4210 -24
rect 33 -57 3437 -40
rect 33 -73 1776 -57
rect 33 -90 971 -73
rect 33 -286 214 -90
rect 433 -269 971 -90
rect 1190 -253 1776 -73
rect 1995 -253 2697 -57
rect 2916 -236 3437 -57
rect 3656 -220 4210 -40
rect 4429 -204 4933 -24
rect 5152 -204 5607 -8
rect 5826 -24 6840 -8
rect 5826 -204 6265 -24
rect 4429 -220 6265 -204
rect 6484 -220 6840 -24
rect 3656 -236 6840 -220
rect 2916 -253 6840 -236
rect 1190 -269 6840 -253
rect 433 -286 6840 -269
rect 33 -1075 6840 -286
<< via3 >>
rect 280 7248 376 7349
rect 539 7248 635 7349
rect 801 7248 897 7349
rect 1048 7251 1144 7352
rect 1300 7252 1396 7353
rect 1552 7251 1648 7352
rect 1801 7251 1897 7352
rect 4400 7261 4496 7362
rect 4743 7261 4839 7362
rect 5098 7273 5194 7374
rect 5398 7277 5494 7378
rect 5613 7285 5709 7386
rect 5890 7261 5986 7362
rect 6088 7300 6184 7401
rect 6272 7288 6368 7389
rect -327 5897 -231 5998
rect -327 5104 -231 5205
rect 7136 6128 7232 6229
rect 7128 5851 7224 5952
rect 7120 5542 7216 5643
rect 7120 5257 7216 5358
rect 7104 5019 7200 5120
rect 7120 4893 7216 4994
rect -343 4294 -247 4395
rect -310 3649 -214 3750
rect -310 3186 -214 3287
rect -294 2674 -198 2775
rect -310 2161 -214 2262
rect -310 1682 -214 1783
rect -277 1202 -181 1303
rect -310 690 -214 791
rect 7076 2240 7295 2436
rect 7072 1865 7291 2061
rect 7080 1497 7299 1693
rect 7084 1221 7303 1417
rect 7092 977 7311 1173
rect 214 -286 433 -90
rect 971 -269 1190 -73
rect 1776 -253 1995 -57
rect 2697 -253 2916 -57
rect 3437 -236 3656 -40
rect 4210 -220 4429 -24
rect 4933 -204 5152 -8
rect 5607 -204 5826 -8
rect 6265 -220 6484 -24
<< metal4 >>
rect 100 7353 2205 7990
rect 100 7352 1300 7353
rect 100 7349 1048 7352
rect 100 7248 280 7349
rect 376 7248 539 7349
rect 635 7248 801 7349
rect 897 7251 1048 7349
rect 1144 7252 1300 7352
rect 1396 7352 2205 7353
rect 1396 7252 1552 7352
rect 1144 7251 1552 7252
rect 1648 7251 1801 7352
rect 1897 7251 2205 7352
rect 897 7248 2205 7251
rect 100 7147 2205 7248
rect 4262 7401 6571 7890
rect 4262 7386 6088 7401
rect 4262 7378 5613 7386
rect 4262 7374 5398 7378
rect 4262 7362 5098 7374
rect 4262 7261 4400 7362
rect 4496 7261 4743 7362
rect 4839 7273 5098 7362
rect 5194 7277 5398 7374
rect 5494 7285 5613 7378
rect 5709 7362 6088 7386
rect 5709 7285 5890 7362
rect 5494 7277 5890 7285
rect 5194 7273 5890 7277
rect 4839 7261 5890 7273
rect 5986 7300 6088 7362
rect 6184 7389 6571 7401
rect 6184 7300 6272 7389
rect 5986 7288 6272 7300
rect 6368 7288 6571 7389
rect 5986 7261 6571 7288
rect 4262 7227 6571 7261
rect -1348 5998 -145 6344
rect -1348 5897 -327 5998
rect -231 5897 -145 5998
rect -1348 5205 -145 5897
rect -1348 5104 -327 5205
rect -231 5104 -145 5205
rect -1348 4395 -145 5104
rect 7080 6229 8221 6319
rect 7080 6128 7136 6229
rect 7232 6128 8221 6229
rect 7080 5952 8221 6128
rect 7080 5851 7128 5952
rect 7224 5851 8221 5952
rect 7080 5643 8221 5851
rect 7080 5542 7120 5643
rect 7216 5542 8221 5643
rect 7080 5358 8221 5542
rect 7080 5257 7120 5358
rect 7216 5257 8221 5358
rect 7080 5120 8221 5257
rect 7080 5019 7104 5120
rect 7200 5019 8221 5120
rect 7080 4994 8221 5019
rect 7080 4893 7120 4994
rect 7216 4893 8221 4994
rect 7080 4718 8221 4893
rect -1348 4294 -343 4395
rect -247 4294 -145 4395
rect -1348 3750 -145 4294
rect -1348 3649 -310 3750
rect -214 3649 -145 3750
rect -1348 3287 -145 3649
rect -1348 3186 -310 3287
rect -214 3186 -145 3287
rect -1348 2775 -145 3186
rect -1348 2674 -294 2775
rect -198 2674 -145 2775
rect -1348 2262 -145 2674
rect -1348 2161 -310 2262
rect -214 2161 -145 2262
rect -1348 1783 -145 2161
rect -1348 1682 -310 1783
rect -214 1682 -145 1783
rect -1348 1303 -145 1682
rect -1348 1202 -277 1303
rect -181 1202 -145 1303
rect -1348 791 -145 1202
rect -1348 690 -310 791
rect -214 690 -145 791
rect 7048 2436 7915 2464
rect 7048 2240 7076 2436
rect 7295 2240 7915 2436
rect 7048 2061 7915 2240
rect 7048 1865 7072 2061
rect 7291 1865 7915 2061
rect 7048 1693 7915 1865
rect 7048 1497 7080 1693
rect 7299 1497 7915 1693
rect 7048 1417 7915 1497
rect 7048 1221 7084 1417
rect 7303 1221 7915 1417
rect 7048 1173 7915 1221
rect 7048 977 7092 1173
rect 7311 977 7915 1173
rect 7048 737 7915 977
rect -1348 339 -145 690
rect 33 -8 6840 158
rect 33 -24 4933 -8
rect 33 -40 4210 -24
rect 33 -57 3437 -40
rect 33 -73 1776 -57
rect 33 -90 971 -73
rect 33 -286 214 -90
rect 433 -269 971 -90
rect 1190 -253 1776 -73
rect 1995 -253 2697 -57
rect 2916 -236 3437 -57
rect 3656 -220 4210 -40
rect 4429 -204 4933 -24
rect 5152 -204 5607 -8
rect 5826 -24 6840 -8
rect 5826 -204 6265 -24
rect 4429 -220 6265 -204
rect 6484 -220 6840 -24
rect 3656 -236 6840 -220
rect 2916 -253 6840 -236
rect 1190 -269 6840 -253
rect 433 -286 6840 -269
rect 33 -1075 6840 -286
use BGR  BGR_0
timestamp 1635312588
transform 1 0 2634 0 1 4394
box -2634 -4394 4277 2732
<< end >>
