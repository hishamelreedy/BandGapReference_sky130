magic
tech sky130A
magscale 1 2
timestamp 1634672276
<< nwell >>
rect 2846 256 2950 388
<< metal1 >>
rect -1294 946 -980 956
rect -1294 932 3018 946
rect -3774 762 3018 932
rect -3774 758 -980 762
rect -3774 328 -3402 758
rect -3774 -3168 -3406 328
rect -3774 -3458 -2540 -3168
<< metal2 >>
rect -5144 4972 8554 5464
rect 2428 3860 2692 4972
rect 3494 3886 3758 4972
rect 4322 3886 4586 4972
rect 5024 3886 5288 4972
rect 4758 412 6192 418
rect 2836 240 2952 396
rect 3000 344 3108 394
rect 3000 258 3022 344
rect 3090 258 3108 344
rect 2868 -108 2932 240
rect 3000 226 3108 258
rect 3776 206 3892 234
rect 3776 120 3798 206
rect 3866 120 3892 206
rect 3776 78 3892 120
rect 3998 180 4092 242
rect 4758 230 6198 412
rect 3998 174 4684 180
rect 3998 76 4804 174
rect 2868 -184 3466 -108
rect 3286 -634 3460 -184
rect 4548 -754 4804 76
rect 5902 -844 6198 230
rect -274 -8274 -136 -6058
rect -5238 -8766 8460 -8274
<< via2 >>
rect 3442 970 3510 1056
rect 3022 258 3090 344
rect 3798 120 3866 206
rect 2020 -932 2088 -846
rect 6936 -984 7004 -898
rect 592 -1474 660 -1388
<< metal3 >>
rect 3428 1056 7090 1074
rect 3428 970 3442 1056
rect 3510 970 7090 1056
rect 3428 940 7090 970
rect 3002 344 3106 358
rect 3002 258 3022 344
rect 3090 258 3106 344
rect 3002 234 3106 258
rect 3014 176 3088 234
rect 3786 206 3880 224
rect 3014 172 3086 176
rect 1992 -268 2900 -264
rect 3016 -268 3086 172
rect 3786 120 3798 206
rect 3866 120 3880 206
rect 3786 112 3880 120
rect 3786 92 3882 112
rect 3790 6 3882 92
rect 1992 -328 3086 -268
rect 1992 -332 3084 -328
rect 1992 -846 2118 -332
rect 1992 -932 2020 -846
rect 2088 -932 2118 -846
rect 1992 -978 2118 -932
rect 3792 -1316 3882 6
rect 6898 -898 7090 940
rect 6898 -984 6936 -898
rect 7004 -984 7090 -898
rect 6898 -1028 7090 -984
rect 530 -1388 3884 -1316
rect 530 -1474 592 -1388
rect 660 -1474 3884 -1388
rect 530 -1538 3884 -1474
use pmos_mirror  pmos_mirror_0
timestamp 1634671827
transform 1 0 4180 0 1 2174
box -4180 -2174 3034 2473
use PDN  PDN_0
timestamp 1634672276
transform 1 0 6158 0 1 -4980
box -11370 -3742 1046 4526
<< labels >>
flabel metal2 -5144 4972 8554 5464 0 FreeSans 1600 0 0 0 VDD!
flabel metal2 -5238 -8766 8460 -8274 0 FreeSans 1600 0 0 0 GND!
<< end >>
