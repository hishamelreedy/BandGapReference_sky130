magic
tech sky130A
magscale 1 2
timestamp 1629311173
<< checkpaint >>
rect -1260 -1260 1956 2474
<< nwell >>
rect 0 0 696 1214
<< pmos >>
rect 204 102 234 1112
rect 290 102 320 1112
rect 376 102 406 1112
rect 462 102 492 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 234 1100 290 1112
rect 234 1066 245 1100
rect 279 1066 290 1100
rect 234 1032 290 1066
rect 234 998 245 1032
rect 279 998 290 1032
rect 234 964 290 998
rect 234 930 245 964
rect 279 930 290 964
rect 234 896 290 930
rect 234 862 245 896
rect 279 862 290 896
rect 234 828 290 862
rect 234 794 245 828
rect 279 794 290 828
rect 234 760 290 794
rect 234 726 245 760
rect 279 726 290 760
rect 234 692 290 726
rect 234 658 245 692
rect 279 658 290 692
rect 234 624 290 658
rect 234 590 245 624
rect 279 590 290 624
rect 234 556 290 590
rect 234 522 245 556
rect 279 522 290 556
rect 234 488 290 522
rect 234 454 245 488
rect 279 454 290 488
rect 234 420 290 454
rect 234 386 245 420
rect 279 386 290 420
rect 234 352 290 386
rect 234 318 245 352
rect 279 318 290 352
rect 234 284 290 318
rect 234 250 245 284
rect 279 250 290 284
rect 234 216 290 250
rect 234 182 245 216
rect 279 182 290 216
rect 234 148 290 182
rect 234 114 245 148
rect 279 114 290 148
rect 234 102 290 114
rect 320 1100 376 1112
rect 320 1066 331 1100
rect 365 1066 376 1100
rect 320 1032 376 1066
rect 320 998 331 1032
rect 365 998 376 1032
rect 320 964 376 998
rect 320 930 331 964
rect 365 930 376 964
rect 320 896 376 930
rect 320 862 331 896
rect 365 862 376 896
rect 320 828 376 862
rect 320 794 331 828
rect 365 794 376 828
rect 320 760 376 794
rect 320 726 331 760
rect 365 726 376 760
rect 320 692 376 726
rect 320 658 331 692
rect 365 658 376 692
rect 320 624 376 658
rect 320 590 331 624
rect 365 590 376 624
rect 320 556 376 590
rect 320 522 331 556
rect 365 522 376 556
rect 320 488 376 522
rect 320 454 331 488
rect 365 454 376 488
rect 320 420 376 454
rect 320 386 331 420
rect 365 386 376 420
rect 320 352 376 386
rect 320 318 331 352
rect 365 318 376 352
rect 320 284 376 318
rect 320 250 331 284
rect 365 250 376 284
rect 320 216 376 250
rect 320 182 331 216
rect 365 182 376 216
rect 320 148 376 182
rect 320 114 331 148
rect 365 114 376 148
rect 320 102 376 114
rect 406 1100 462 1112
rect 406 1066 417 1100
rect 451 1066 462 1100
rect 406 1032 462 1066
rect 406 998 417 1032
rect 451 998 462 1032
rect 406 964 462 998
rect 406 930 417 964
rect 451 930 462 964
rect 406 896 462 930
rect 406 862 417 896
rect 451 862 462 896
rect 406 828 462 862
rect 406 794 417 828
rect 451 794 462 828
rect 406 760 462 794
rect 406 726 417 760
rect 451 726 462 760
rect 406 692 462 726
rect 406 658 417 692
rect 451 658 462 692
rect 406 624 462 658
rect 406 590 417 624
rect 451 590 462 624
rect 406 556 462 590
rect 406 522 417 556
rect 451 522 462 556
rect 406 488 462 522
rect 406 454 417 488
rect 451 454 462 488
rect 406 420 462 454
rect 406 386 417 420
rect 451 386 462 420
rect 406 352 462 386
rect 406 318 417 352
rect 451 318 462 352
rect 406 284 462 318
rect 406 250 417 284
rect 451 250 462 284
rect 406 216 462 250
rect 406 182 417 216
rect 451 182 462 216
rect 406 148 462 182
rect 406 114 417 148
rect 451 114 462 148
rect 406 102 462 114
rect 492 1100 548 1112
rect 492 1066 503 1100
rect 537 1066 548 1100
rect 492 1032 548 1066
rect 492 998 503 1032
rect 537 998 548 1032
rect 492 964 548 998
rect 492 930 503 964
rect 537 930 548 964
rect 492 896 548 930
rect 492 862 503 896
rect 537 862 548 896
rect 492 828 548 862
rect 492 794 503 828
rect 537 794 548 828
rect 492 760 548 794
rect 492 726 503 760
rect 537 726 548 760
rect 492 692 548 726
rect 492 658 503 692
rect 537 658 548 692
rect 492 624 548 658
rect 492 590 503 624
rect 537 590 548 624
rect 492 556 548 590
rect 492 522 503 556
rect 537 522 548 556
rect 492 488 548 522
rect 492 454 503 488
rect 537 454 548 488
rect 492 420 548 454
rect 492 386 503 420
rect 537 386 548 420
rect 492 352 548 386
rect 492 318 503 352
rect 537 318 548 352
rect 492 284 548 318
rect 492 250 503 284
rect 537 250 548 284
rect 492 216 548 250
rect 492 182 503 216
rect 537 182 548 216
rect 492 148 548 182
rect 492 114 503 148
rect 537 114 548 148
rect 492 102 548 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 245 1066 279 1100
rect 245 998 279 1032
rect 245 930 279 964
rect 245 862 279 896
rect 245 794 279 828
rect 245 726 279 760
rect 245 658 279 692
rect 245 590 279 624
rect 245 522 279 556
rect 245 454 279 488
rect 245 386 279 420
rect 245 318 279 352
rect 245 250 279 284
rect 245 182 279 216
rect 245 114 279 148
rect 331 1066 365 1100
rect 331 998 365 1032
rect 331 930 365 964
rect 331 862 365 896
rect 331 794 365 828
rect 331 726 365 760
rect 331 658 365 692
rect 331 590 365 624
rect 331 522 365 556
rect 331 454 365 488
rect 331 386 365 420
rect 331 318 365 352
rect 331 250 365 284
rect 331 182 365 216
rect 331 114 365 148
rect 417 1066 451 1100
rect 417 998 451 1032
rect 417 930 451 964
rect 417 862 451 896
rect 417 794 451 828
rect 417 726 451 760
rect 417 658 451 692
rect 417 590 451 624
rect 417 522 451 556
rect 417 454 451 488
rect 417 386 451 420
rect 417 318 451 352
rect 417 250 451 284
rect 417 182 451 216
rect 417 114 451 148
rect 503 1066 537 1100
rect 503 998 537 1032
rect 503 930 537 964
rect 503 862 537 896
rect 503 794 537 828
rect 503 726 537 760
rect 503 658 537 692
rect 503 590 537 624
rect 503 522 537 556
rect 503 454 537 488
rect 503 386 537 420
rect 503 318 537 352
rect 503 250 537 284
rect 503 182 537 216
rect 503 114 537 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 602 1066 660 1112
rect 602 1032 614 1066
rect 648 1032 660 1066
rect 602 998 660 1032
rect 602 964 614 998
rect 648 964 660 998
rect 602 930 660 964
rect 602 896 614 930
rect 648 896 660 930
rect 602 862 660 896
rect 602 828 614 862
rect 648 828 660 862
rect 602 794 660 828
rect 602 760 614 794
rect 648 760 660 794
rect 602 726 660 760
rect 602 692 614 726
rect 648 692 660 726
rect 602 658 660 692
rect 602 624 614 658
rect 648 624 660 658
rect 602 590 660 624
rect 602 556 614 590
rect 648 556 660 590
rect 602 522 660 556
rect 602 488 614 522
rect 648 488 660 522
rect 602 454 660 488
rect 602 420 614 454
rect 648 420 660 454
rect 602 386 660 420
rect 602 352 614 386
rect 648 352 660 386
rect 602 318 660 352
rect 602 284 614 318
rect 648 284 660 318
rect 602 250 660 284
rect 602 216 614 250
rect 648 216 660 250
rect 602 182 660 216
rect 602 148 614 182
rect 648 148 660 182
rect 602 102 660 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 614 1032 648 1066
rect 614 964 648 998
rect 614 896 648 930
rect 614 828 648 862
rect 614 760 648 794
rect 614 692 648 726
rect 614 624 648 658
rect 614 556 648 590
rect 614 488 648 522
rect 614 420 648 454
rect 614 352 648 386
rect 614 284 648 318
rect 614 216 648 250
rect 614 148 648 182
<< poly >>
rect 179 1194 517 1214
rect 179 1160 195 1194
rect 229 1160 263 1194
rect 297 1160 331 1194
rect 365 1160 399 1194
rect 433 1160 467 1194
rect 501 1160 517 1194
rect 179 1144 517 1160
rect 204 1112 234 1144
rect 290 1112 320 1144
rect 376 1112 406 1144
rect 462 1112 492 1144
rect 204 70 234 102
rect 290 70 320 102
rect 376 70 406 102
rect 462 70 492 102
rect 179 54 517 70
rect 179 20 195 54
rect 229 20 263 54
rect 297 20 331 54
rect 365 20 399 54
rect 433 20 467 54
rect 501 20 517 54
rect 179 0 517 20
<< polycont >>
rect 195 1160 229 1194
rect 263 1160 297 1194
rect 331 1160 365 1194
rect 399 1160 433 1194
rect 467 1160 501 1194
rect 195 20 229 54
rect 263 20 297 54
rect 331 20 365 54
rect 399 20 433 54
rect 467 20 501 54
<< locali >>
rect 179 1160 187 1194
rect 229 1160 259 1194
rect 297 1160 331 1194
rect 365 1160 399 1194
rect 437 1160 467 1194
rect 509 1160 517 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 245 1100 279 1116
rect 245 1032 279 1058
rect 245 964 279 986
rect 245 896 279 914
rect 245 828 279 842
rect 245 760 279 770
rect 245 692 279 698
rect 245 624 279 626
rect 245 588 279 590
rect 245 516 279 522
rect 245 444 279 454
rect 245 372 279 386
rect 245 300 279 318
rect 245 228 279 250
rect 245 156 279 182
rect 245 98 279 114
rect 331 1100 365 1116
rect 331 1032 365 1058
rect 331 964 365 986
rect 331 896 365 914
rect 331 828 365 842
rect 331 760 365 770
rect 331 692 365 698
rect 331 624 365 626
rect 331 588 365 590
rect 331 516 365 522
rect 331 444 365 454
rect 331 372 365 386
rect 331 300 365 318
rect 331 228 365 250
rect 331 156 365 182
rect 331 98 365 114
rect 417 1100 451 1116
rect 417 1032 451 1058
rect 417 964 451 986
rect 417 896 451 914
rect 417 828 451 842
rect 417 760 451 770
rect 417 692 451 698
rect 417 624 451 626
rect 417 588 451 590
rect 417 516 451 522
rect 417 444 451 454
rect 417 372 451 386
rect 417 300 451 318
rect 417 228 451 250
rect 417 156 451 182
rect 417 98 451 114
rect 503 1100 537 1116
rect 503 1032 537 1058
rect 503 964 537 986
rect 503 896 537 914
rect 503 828 537 842
rect 503 760 537 770
rect 503 692 537 698
rect 503 624 537 626
rect 503 588 537 590
rect 503 516 537 522
rect 503 444 537 454
rect 503 372 537 386
rect 503 300 537 318
rect 503 228 537 250
rect 503 156 537 182
rect 614 1020 648 1032
rect 614 948 648 964
rect 614 876 648 896
rect 614 804 648 828
rect 614 732 648 760
rect 614 660 648 692
rect 614 590 648 624
rect 614 522 648 554
rect 614 454 648 482
rect 614 386 648 410
rect 614 318 648 338
rect 614 250 648 266
rect 614 182 648 194
rect 503 98 537 114
rect 179 20 187 54
rect 229 20 259 54
rect 297 20 331 54
rect 365 20 399 54
rect 437 20 467 54
rect 509 20 517 54
<< viali >>
rect 187 1160 195 1194
rect 195 1160 221 1194
rect 259 1160 263 1194
rect 263 1160 293 1194
rect 331 1160 365 1194
rect 403 1160 433 1194
rect 433 1160 437 1194
rect 475 1160 501 1194
rect 501 1160 509 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 245 1066 279 1092
rect 245 1058 279 1066
rect 245 998 279 1020
rect 245 986 279 998
rect 245 930 279 948
rect 245 914 279 930
rect 245 862 279 876
rect 245 842 279 862
rect 245 794 279 804
rect 245 770 279 794
rect 245 726 279 732
rect 245 698 279 726
rect 245 658 279 660
rect 245 626 279 658
rect 245 556 279 588
rect 245 554 279 556
rect 245 488 279 516
rect 245 482 279 488
rect 245 420 279 444
rect 245 410 279 420
rect 245 352 279 372
rect 245 338 279 352
rect 245 284 279 300
rect 245 266 279 284
rect 245 216 279 228
rect 245 194 279 216
rect 245 148 279 156
rect 245 122 279 148
rect 331 1066 365 1092
rect 331 1058 365 1066
rect 331 998 365 1020
rect 331 986 365 998
rect 331 930 365 948
rect 331 914 365 930
rect 331 862 365 876
rect 331 842 365 862
rect 331 794 365 804
rect 331 770 365 794
rect 331 726 365 732
rect 331 698 365 726
rect 331 658 365 660
rect 331 626 365 658
rect 331 556 365 588
rect 331 554 365 556
rect 331 488 365 516
rect 331 482 365 488
rect 331 420 365 444
rect 331 410 365 420
rect 331 352 365 372
rect 331 338 365 352
rect 331 284 365 300
rect 331 266 365 284
rect 331 216 365 228
rect 331 194 365 216
rect 331 148 365 156
rect 331 122 365 148
rect 417 1066 451 1092
rect 417 1058 451 1066
rect 417 998 451 1020
rect 417 986 451 998
rect 417 930 451 948
rect 417 914 451 930
rect 417 862 451 876
rect 417 842 451 862
rect 417 794 451 804
rect 417 770 451 794
rect 417 726 451 732
rect 417 698 451 726
rect 417 658 451 660
rect 417 626 451 658
rect 417 556 451 588
rect 417 554 451 556
rect 417 488 451 516
rect 417 482 451 488
rect 417 420 451 444
rect 417 410 451 420
rect 417 352 451 372
rect 417 338 451 352
rect 417 284 451 300
rect 417 266 451 284
rect 417 216 451 228
rect 417 194 451 216
rect 417 148 451 156
rect 417 122 451 148
rect 503 1066 537 1092
rect 503 1058 537 1066
rect 503 998 537 1020
rect 503 986 537 998
rect 503 930 537 948
rect 503 914 537 930
rect 503 862 537 876
rect 503 842 537 862
rect 503 794 537 804
rect 503 770 537 794
rect 503 726 537 732
rect 503 698 537 726
rect 503 658 537 660
rect 503 626 537 658
rect 503 556 537 588
rect 503 554 537 556
rect 503 488 537 516
rect 503 482 537 488
rect 503 420 537 444
rect 503 410 537 420
rect 503 352 537 372
rect 503 338 537 352
rect 503 284 537 300
rect 503 266 537 284
rect 503 216 537 228
rect 503 194 537 216
rect 503 148 537 156
rect 503 122 537 148
rect 614 1066 648 1092
rect 614 1058 648 1066
rect 614 998 648 1020
rect 614 986 648 998
rect 614 930 648 948
rect 614 914 648 930
rect 614 862 648 876
rect 614 842 648 862
rect 614 794 648 804
rect 614 770 648 794
rect 614 726 648 732
rect 614 698 648 726
rect 614 658 648 660
rect 614 626 648 658
rect 614 556 648 588
rect 614 554 648 556
rect 614 488 648 516
rect 614 482 648 488
rect 614 420 648 444
rect 614 410 648 420
rect 614 352 648 372
rect 614 338 648 352
rect 614 284 648 300
rect 614 266 648 284
rect 614 216 648 228
rect 614 194 648 216
rect 614 148 648 156
rect 614 122 648 148
rect 187 20 195 54
rect 195 20 221 54
rect 259 20 263 54
rect 263 20 293 54
rect 331 20 365 54
rect 403 20 433 54
rect 433 20 437 54
rect 475 20 501 54
rect 501 20 509 54
<< metal1 >>
rect 175 1194 521 1214
rect 175 1160 187 1194
rect 221 1160 259 1194
rect 293 1160 331 1194
rect 365 1160 403 1194
rect 437 1160 475 1194
rect 509 1160 521 1194
rect 175 1148 521 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 236 1098 288 1104
rect 236 1034 288 1046
rect 236 970 288 982
rect 236 914 245 918
rect 279 914 288 918
rect 236 906 288 914
rect 236 842 245 854
rect 279 842 288 854
rect 236 778 245 790
rect 279 778 288 790
rect 236 714 245 726
rect 279 714 288 726
rect 236 660 288 662
rect 236 626 245 660
rect 279 626 288 660
rect 236 588 288 626
rect 236 554 245 588
rect 279 554 288 588
rect 236 516 288 554
rect 236 482 245 516
rect 279 482 288 516
rect 236 444 288 482
rect 236 410 245 444
rect 279 410 288 444
rect 236 372 288 410
rect 236 338 245 372
rect 279 338 288 372
rect 236 300 288 338
rect 236 266 245 300
rect 279 266 288 300
rect 236 228 288 266
rect 236 194 245 228
rect 279 194 288 228
rect 236 156 288 194
rect 236 122 245 156
rect 279 122 288 156
rect 236 110 288 122
rect 322 1092 374 1104
rect 322 1058 331 1092
rect 365 1058 374 1092
rect 322 1020 374 1058
rect 322 986 331 1020
rect 365 986 374 1020
rect 322 948 374 986
rect 322 914 331 948
rect 365 914 374 948
rect 322 876 374 914
rect 322 842 331 876
rect 365 842 374 876
rect 322 804 374 842
rect 322 770 331 804
rect 365 770 374 804
rect 322 732 374 770
rect 322 698 331 732
rect 365 698 374 732
rect 322 660 374 698
rect 322 626 331 660
rect 365 626 374 660
rect 322 588 374 626
rect 322 554 331 588
rect 365 554 374 588
rect 322 552 374 554
rect 322 488 331 500
rect 365 488 374 500
rect 322 424 331 436
rect 365 424 374 436
rect 322 360 331 372
rect 365 360 374 372
rect 322 300 374 308
rect 322 296 331 300
rect 365 296 374 300
rect 322 232 374 244
rect 322 168 374 180
rect 322 110 374 116
rect 408 1098 460 1104
rect 408 1034 460 1046
rect 408 970 460 982
rect 408 914 417 918
rect 451 914 460 918
rect 408 906 460 914
rect 408 842 417 854
rect 451 842 460 854
rect 408 778 417 790
rect 451 778 460 790
rect 408 714 417 726
rect 451 714 460 726
rect 408 660 460 662
rect 408 626 417 660
rect 451 626 460 660
rect 408 588 460 626
rect 408 554 417 588
rect 451 554 460 588
rect 408 516 460 554
rect 408 482 417 516
rect 451 482 460 516
rect 408 444 460 482
rect 408 410 417 444
rect 451 410 460 444
rect 408 372 460 410
rect 408 338 417 372
rect 451 338 460 372
rect 408 300 460 338
rect 408 266 417 300
rect 451 266 460 300
rect 408 228 460 266
rect 408 194 417 228
rect 451 194 460 228
rect 408 156 460 194
rect 408 122 417 156
rect 451 122 460 156
rect 408 110 460 122
rect 494 1092 546 1104
rect 494 1058 503 1092
rect 537 1058 546 1092
rect 494 1020 546 1058
rect 494 986 503 1020
rect 537 986 546 1020
rect 494 948 546 986
rect 494 914 503 948
rect 537 914 546 948
rect 494 876 546 914
rect 494 842 503 876
rect 537 842 546 876
rect 494 804 546 842
rect 494 770 503 804
rect 537 770 546 804
rect 494 732 546 770
rect 494 698 503 732
rect 537 698 546 732
rect 494 660 546 698
rect 494 626 503 660
rect 537 626 546 660
rect 494 588 546 626
rect 494 554 503 588
rect 537 554 546 588
rect 494 552 546 554
rect 494 488 503 500
rect 537 488 546 500
rect 494 424 503 436
rect 537 424 546 436
rect 494 360 503 372
rect 537 360 546 372
rect 494 300 546 308
rect 494 296 503 300
rect 537 296 546 300
rect 494 232 546 244
rect 494 168 546 180
rect 494 110 546 116
rect 602 1092 660 1104
rect 602 1058 614 1092
rect 648 1058 660 1092
rect 602 1020 660 1058
rect 602 986 614 1020
rect 648 986 660 1020
rect 602 948 660 986
rect 602 914 614 948
rect 648 914 660 948
rect 602 876 660 914
rect 602 842 614 876
rect 648 842 660 876
rect 602 804 660 842
rect 602 770 614 804
rect 648 770 660 804
rect 602 732 660 770
rect 602 698 614 732
rect 648 698 660 732
rect 602 660 660 698
rect 602 626 614 660
rect 648 626 660 660
rect 602 588 660 626
rect 602 554 614 588
rect 648 554 660 588
rect 602 516 660 554
rect 602 482 614 516
rect 648 482 660 516
rect 602 444 660 482
rect 602 410 614 444
rect 648 410 660 444
rect 602 372 660 410
rect 602 338 614 372
rect 648 338 660 372
rect 602 300 660 338
rect 602 266 614 300
rect 648 266 660 300
rect 602 228 660 266
rect 602 194 614 228
rect 648 194 660 228
rect 602 156 660 194
rect 602 122 614 156
rect 648 122 660 156
rect 602 110 660 122
rect 175 54 521 66
rect 175 20 187 54
rect 221 20 259 54
rect 293 20 331 54
rect 365 20 403 54
rect 437 20 475 54
rect 509 20 521 54
rect 175 0 521 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 236 1092 288 1098
rect 236 1058 245 1092
rect 245 1058 279 1092
rect 279 1058 288 1092
rect 236 1046 288 1058
rect 236 1020 288 1034
rect 236 986 245 1020
rect 245 986 279 1020
rect 279 986 288 1020
rect 236 982 288 986
rect 236 948 288 970
rect 236 918 245 948
rect 245 918 279 948
rect 279 918 288 948
rect 236 876 288 906
rect 236 854 245 876
rect 245 854 279 876
rect 279 854 288 876
rect 236 804 288 842
rect 236 790 245 804
rect 245 790 279 804
rect 279 790 288 804
rect 236 770 245 778
rect 245 770 279 778
rect 279 770 288 778
rect 236 732 288 770
rect 236 726 245 732
rect 245 726 279 732
rect 279 726 288 732
rect 236 698 245 714
rect 245 698 279 714
rect 279 698 288 714
rect 236 662 288 698
rect 322 516 374 552
rect 322 500 331 516
rect 331 500 365 516
rect 365 500 374 516
rect 322 482 331 488
rect 331 482 365 488
rect 365 482 374 488
rect 322 444 374 482
rect 322 436 331 444
rect 331 436 365 444
rect 365 436 374 444
rect 322 410 331 424
rect 331 410 365 424
rect 365 410 374 424
rect 322 372 374 410
rect 322 338 331 360
rect 331 338 365 360
rect 365 338 374 360
rect 322 308 374 338
rect 322 266 331 296
rect 331 266 365 296
rect 365 266 374 296
rect 322 244 374 266
rect 322 228 374 232
rect 322 194 331 228
rect 331 194 365 228
rect 365 194 374 228
rect 322 180 374 194
rect 322 156 374 168
rect 322 122 331 156
rect 331 122 365 156
rect 365 122 374 156
rect 322 116 374 122
rect 408 1092 460 1098
rect 408 1058 417 1092
rect 417 1058 451 1092
rect 451 1058 460 1092
rect 408 1046 460 1058
rect 408 1020 460 1034
rect 408 986 417 1020
rect 417 986 451 1020
rect 451 986 460 1020
rect 408 982 460 986
rect 408 948 460 970
rect 408 918 417 948
rect 417 918 451 948
rect 451 918 460 948
rect 408 876 460 906
rect 408 854 417 876
rect 417 854 451 876
rect 451 854 460 876
rect 408 804 460 842
rect 408 790 417 804
rect 417 790 451 804
rect 451 790 460 804
rect 408 770 417 778
rect 417 770 451 778
rect 451 770 460 778
rect 408 732 460 770
rect 408 726 417 732
rect 417 726 451 732
rect 451 726 460 732
rect 408 698 417 714
rect 417 698 451 714
rect 451 698 460 714
rect 408 662 460 698
rect 494 516 546 552
rect 494 500 503 516
rect 503 500 537 516
rect 537 500 546 516
rect 494 482 503 488
rect 503 482 537 488
rect 537 482 546 488
rect 494 444 546 482
rect 494 436 503 444
rect 503 436 537 444
rect 537 436 546 444
rect 494 410 503 424
rect 503 410 537 424
rect 537 410 546 424
rect 494 372 546 410
rect 494 338 503 360
rect 503 338 537 360
rect 537 338 546 360
rect 494 308 546 338
rect 494 266 503 296
rect 503 266 537 296
rect 537 266 546 296
rect 494 244 546 266
rect 494 228 546 232
rect 494 194 503 228
rect 503 194 537 228
rect 537 194 546 228
rect 494 180 546 194
rect 494 156 546 168
rect 494 122 503 156
rect 503 122 537 156
rect 537 122 546 156
rect 494 116 546 122
<< metal2 >>
rect 10 1098 686 1104
rect 10 1046 236 1098
rect 288 1046 408 1098
rect 460 1046 686 1098
rect 10 1034 686 1046
rect 10 982 236 1034
rect 288 982 408 1034
rect 460 982 686 1034
rect 10 970 686 982
rect 10 918 236 970
rect 288 918 408 970
rect 460 918 686 970
rect 10 906 686 918
rect 10 854 236 906
rect 288 854 408 906
rect 460 854 686 906
rect 10 842 686 854
rect 10 790 236 842
rect 288 790 408 842
rect 460 790 686 842
rect 10 778 686 790
rect 10 726 236 778
rect 288 726 408 778
rect 460 726 686 778
rect 10 714 686 726
rect 10 662 236 714
rect 288 662 408 714
rect 460 662 686 714
rect 10 632 686 662
rect 10 552 686 582
rect 10 500 150 552
rect 202 500 322 552
rect 374 500 494 552
rect 546 500 686 552
rect 10 488 686 500
rect 10 436 150 488
rect 202 436 322 488
rect 374 436 494 488
rect 546 436 686 488
rect 10 424 686 436
rect 10 372 150 424
rect 202 372 322 424
rect 374 372 494 424
rect 546 372 686 424
rect 10 360 686 372
rect 10 308 150 360
rect 202 308 322 360
rect 374 308 494 360
rect 546 308 686 360
rect 10 296 686 308
rect 10 244 150 296
rect 202 244 322 296
rect 374 244 494 296
rect 546 244 686 296
rect 10 232 686 244
rect 10 180 150 232
rect 202 180 322 232
rect 374 180 494 232
rect 546 180 686 232
rect 10 168 686 180
rect 10 116 150 168
rect 202 116 322 168
rect 374 116 494 168
rect 546 116 686 168
rect 10 110 686 116
<< labels >>
flabel comment s 520 607 520 607 0 FreeSans 300 0 0 0 S
flabel comment s 434 607 434 607 0 FreeSans 300 0 0 0 D
flabel comment s 348 607 348 607 0 FreeSans 300 0 0 0 S
flabel comment s 262 607 262 607 0 FreeSans 300 0 0 0 D
flabel comment s 176 607 176 607 0 FreeSans 300 0 0 0 S
flabel comment s 176 607 176 607 0 FreeSans 300 0 0 0 S
flabel comment s 262 607 262 607 0 FreeSans 300 0 0 0 S
flabel comment s 348 607 348 607 0 FreeSans 300 0 0 0 S
flabel comment s 434 607 434 607 0 FreeSans 300 0 0 0 S
flabel metal1 s 326 1170 384 1195 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 330 14 388 39 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 614 605 648 616 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal1 s 48 598 82 609 0 FreeSans 100 0 0 0 BULK
port 1 nsew
flabel metal2 s 60 855 75 921 0 FreeSans 100 0 0 0 DRAIN
port 2 nsew
flabel metal2 s 61 311 75 374 0 FreeSans 100 0 0 0 SOURCE
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9447532
string GDS_START 9425630
<< end >>
