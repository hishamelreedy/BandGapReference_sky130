magic
tech sky130A
magscale 1 2
timestamp 1634505583
<< nwell >>
rect -194 -200 194 200
<< pmoslvt >>
rect -100 -100 100 100
<< pdiff >>
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
<< pdiffc >>
rect -146 -88 -112 88
rect 112 -88 146 88
<< poly >>
rect -58 181 58 197
rect -58 164 -42 181
rect -100 147 -42 164
rect 42 164 58 181
rect 42 147 100 164
rect -100 100 100 147
rect -100 -147 100 -100
rect -100 -164 -42 -147
rect -58 -181 -42 -164
rect 42 -164 100 -147
rect 42 -181 58 -164
rect -58 -197 58 -181
<< polycont >>
rect -42 147 42 181
rect -42 -181 42 -147
<< locali >>
rect -58 147 -42 181
rect 42 147 58 181
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect -58 -181 -42 -147
rect 42 -181 58 -147
<< viali >>
rect -42 147 42 181
rect -146 -88 -112 88
rect 112 -88 146 88
rect -42 -181 42 -147
<< metal1 >>
rect -54 181 54 187
rect -54 147 -42 181
rect 42 147 54 181
rect -54 141 54 147
rect -152 88 -106 100
rect -152 -88 -146 88
rect -112 -88 -106 88
rect -152 -100 -106 -88
rect 106 88 152 100
rect 106 -88 112 88
rect 146 -88 152 88
rect 106 -100 152 -88
rect -54 -147 54 -141
rect -54 -181 -42 -147
rect 42 -181 54 -147
rect -54 -187 54 -181
<< labels >>
flabel pmoslvt -100 -100 100 100 0 FreeSans 800 0 0 0 M9
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 1 l 1 m 1 nf 1 diffcov 100 polycov 50 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
