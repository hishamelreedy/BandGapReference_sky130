magic
tech sky130A
magscale 1 2
timestamp 1622522911
<< nwell >>
rect -2747 -684 2747 684
<< pmoslvt >>
rect -2551 -536 -2351 464
rect -2293 -536 -2093 464
rect -2035 -536 -1835 464
rect -1777 -536 -1577 464
rect -1519 -536 -1319 464
rect -1261 -536 -1061 464
rect -1003 -536 -803 464
rect -745 -536 -545 464
rect -487 -536 -287 464
rect -229 -536 -29 464
rect 29 -536 229 464
rect 287 -536 487 464
rect 545 -536 745 464
rect 803 -536 1003 464
rect 1061 -536 1261 464
rect 1319 -536 1519 464
rect 1577 -536 1777 464
rect 1835 -536 2035 464
rect 2093 -536 2293 464
rect 2351 -536 2551 464
<< pdiff >>
rect -2609 452 -2551 464
rect -2609 -524 -2597 452
rect -2563 -524 -2551 452
rect -2609 -536 -2551 -524
rect -2351 452 -2293 464
rect -2351 -524 -2339 452
rect -2305 -524 -2293 452
rect -2351 -536 -2293 -524
rect -2093 452 -2035 464
rect -2093 -524 -2081 452
rect -2047 -524 -2035 452
rect -2093 -536 -2035 -524
rect -1835 452 -1777 464
rect -1835 -524 -1823 452
rect -1789 -524 -1777 452
rect -1835 -536 -1777 -524
rect -1577 452 -1519 464
rect -1577 -524 -1565 452
rect -1531 -524 -1519 452
rect -1577 -536 -1519 -524
rect -1319 452 -1261 464
rect -1319 -524 -1307 452
rect -1273 -524 -1261 452
rect -1319 -536 -1261 -524
rect -1061 452 -1003 464
rect -1061 -524 -1049 452
rect -1015 -524 -1003 452
rect -1061 -536 -1003 -524
rect -803 452 -745 464
rect -803 -524 -791 452
rect -757 -524 -745 452
rect -803 -536 -745 -524
rect -545 452 -487 464
rect -545 -524 -533 452
rect -499 -524 -487 452
rect -545 -536 -487 -524
rect -287 452 -229 464
rect -287 -524 -275 452
rect -241 -524 -229 452
rect -287 -536 -229 -524
rect -29 452 29 464
rect -29 -524 -17 452
rect 17 -524 29 452
rect -29 -536 29 -524
rect 229 452 287 464
rect 229 -524 241 452
rect 275 -524 287 452
rect 229 -536 287 -524
rect 487 452 545 464
rect 487 -524 499 452
rect 533 -524 545 452
rect 487 -536 545 -524
rect 745 452 803 464
rect 745 -524 757 452
rect 791 -524 803 452
rect 745 -536 803 -524
rect 1003 452 1061 464
rect 1003 -524 1015 452
rect 1049 -524 1061 452
rect 1003 -536 1061 -524
rect 1261 452 1319 464
rect 1261 -524 1273 452
rect 1307 -524 1319 452
rect 1261 -536 1319 -524
rect 1519 452 1577 464
rect 1519 -524 1531 452
rect 1565 -524 1577 452
rect 1519 -536 1577 -524
rect 1777 452 1835 464
rect 1777 -524 1789 452
rect 1823 -524 1835 452
rect 1777 -536 1835 -524
rect 2035 452 2093 464
rect 2035 -524 2047 452
rect 2081 -524 2093 452
rect 2035 -536 2093 -524
rect 2293 452 2351 464
rect 2293 -524 2305 452
rect 2339 -524 2351 452
rect 2293 -536 2351 -524
rect 2551 452 2609 464
rect 2551 -524 2563 452
rect 2597 -524 2609 452
rect 2551 -536 2609 -524
<< pdiffc >>
rect -2597 -524 -2563 452
rect -2339 -524 -2305 452
rect -2081 -524 -2047 452
rect -1823 -524 -1789 452
rect -1565 -524 -1531 452
rect -1307 -524 -1273 452
rect -1049 -524 -1015 452
rect -791 -524 -757 452
rect -533 -524 -499 452
rect -275 -524 -241 452
rect -17 -524 17 452
rect 241 -524 275 452
rect 499 -524 533 452
rect 757 -524 791 452
rect 1015 -524 1049 452
rect 1273 -524 1307 452
rect 1531 -524 1565 452
rect 1789 -524 1823 452
rect 2047 -524 2081 452
rect 2305 -524 2339 452
rect 2563 -524 2597 452
<< nsubdiff >>
rect -2711 614 -2615 648
rect 2615 614 2711 648
rect -2711 551 -2677 614
rect 2677 551 2711 614
rect -2711 -614 -2677 -551
rect 2677 -614 2711 -551
rect -2711 -648 -2615 -614
rect 2615 -648 2711 -614
<< nsubdiffcont >>
rect -2615 614 2615 648
rect -2711 -551 -2677 551
rect 2677 -551 2711 551
rect -2615 -648 2615 -614
<< poly >>
rect -2551 545 -2351 561
rect -2551 511 -2535 545
rect -2367 511 -2351 545
rect -2551 464 -2351 511
rect -2293 545 -2093 561
rect -2293 511 -2277 545
rect -2109 511 -2093 545
rect -2293 464 -2093 511
rect -2035 545 -1835 561
rect -2035 511 -2019 545
rect -1851 511 -1835 545
rect -2035 464 -1835 511
rect -1777 545 -1577 561
rect -1777 511 -1761 545
rect -1593 511 -1577 545
rect -1777 464 -1577 511
rect -1519 545 -1319 561
rect -1519 511 -1503 545
rect -1335 511 -1319 545
rect -1519 464 -1319 511
rect -1261 545 -1061 561
rect -1261 511 -1245 545
rect -1077 511 -1061 545
rect -1261 464 -1061 511
rect -1003 545 -803 561
rect -1003 511 -987 545
rect -819 511 -803 545
rect -1003 464 -803 511
rect -745 545 -545 561
rect -745 511 -729 545
rect -561 511 -545 545
rect -745 464 -545 511
rect -487 545 -287 561
rect -487 511 -471 545
rect -303 511 -287 545
rect -487 464 -287 511
rect -229 545 -29 561
rect -229 511 -213 545
rect -45 511 -29 545
rect -229 464 -29 511
rect 29 545 229 561
rect 29 511 45 545
rect 213 511 229 545
rect 29 464 229 511
rect 287 545 487 561
rect 287 511 303 545
rect 471 511 487 545
rect 287 464 487 511
rect 545 545 745 561
rect 545 511 561 545
rect 729 511 745 545
rect 545 464 745 511
rect 803 545 1003 561
rect 803 511 819 545
rect 987 511 1003 545
rect 803 464 1003 511
rect 1061 545 1261 561
rect 1061 511 1077 545
rect 1245 511 1261 545
rect 1061 464 1261 511
rect 1319 545 1519 561
rect 1319 511 1335 545
rect 1503 511 1519 545
rect 1319 464 1519 511
rect 1577 545 1777 561
rect 1577 511 1593 545
rect 1761 511 1777 545
rect 1577 464 1777 511
rect 1835 545 2035 561
rect 1835 511 1851 545
rect 2019 511 2035 545
rect 1835 464 2035 511
rect 2093 545 2293 561
rect 2093 511 2109 545
rect 2277 511 2293 545
rect 2093 464 2293 511
rect 2351 545 2551 561
rect 2351 511 2367 545
rect 2535 511 2551 545
rect 2351 464 2551 511
rect -2551 -562 -2351 -536
rect -2293 -562 -2093 -536
rect -2035 -562 -1835 -536
rect -1777 -562 -1577 -536
rect -1519 -562 -1319 -536
rect -1261 -562 -1061 -536
rect -1003 -562 -803 -536
rect -745 -562 -545 -536
rect -487 -562 -287 -536
rect -229 -562 -29 -536
rect 29 -562 229 -536
rect 287 -562 487 -536
rect 545 -562 745 -536
rect 803 -562 1003 -536
rect 1061 -562 1261 -536
rect 1319 -562 1519 -536
rect 1577 -562 1777 -536
rect 1835 -562 2035 -536
rect 2093 -562 2293 -536
rect 2351 -562 2551 -536
<< polycont >>
rect -2535 511 -2367 545
rect -2277 511 -2109 545
rect -2019 511 -1851 545
rect -1761 511 -1593 545
rect -1503 511 -1335 545
rect -1245 511 -1077 545
rect -987 511 -819 545
rect -729 511 -561 545
rect -471 511 -303 545
rect -213 511 -45 545
rect 45 511 213 545
rect 303 511 471 545
rect 561 511 729 545
rect 819 511 987 545
rect 1077 511 1245 545
rect 1335 511 1503 545
rect 1593 511 1761 545
rect 1851 511 2019 545
rect 2109 511 2277 545
rect 2367 511 2535 545
<< locali >>
rect -2711 614 -2615 648
rect 2615 614 2711 648
rect -2711 551 -2677 614
rect 2677 551 2711 614
rect -2551 511 -2535 545
rect -2367 511 -2351 545
rect -2293 511 -2277 545
rect -2109 511 -2093 545
rect -2035 511 -2019 545
rect -1851 511 -1835 545
rect -1777 511 -1761 545
rect -1593 511 -1577 545
rect -1519 511 -1503 545
rect -1335 511 -1319 545
rect -1261 511 -1245 545
rect -1077 511 -1061 545
rect -1003 511 -987 545
rect -819 511 -803 545
rect -745 511 -729 545
rect -561 511 -545 545
rect -487 511 -471 545
rect -303 511 -287 545
rect -229 511 -213 545
rect -45 511 -29 545
rect 29 511 45 545
rect 213 511 229 545
rect 287 511 303 545
rect 471 511 487 545
rect 545 511 561 545
rect 729 511 745 545
rect 803 511 819 545
rect 987 511 1003 545
rect 1061 511 1077 545
rect 1245 511 1261 545
rect 1319 511 1335 545
rect 1503 511 1519 545
rect 1577 511 1593 545
rect 1761 511 1777 545
rect 1835 511 1851 545
rect 2019 511 2035 545
rect 2093 511 2109 545
rect 2277 511 2293 545
rect 2351 511 2367 545
rect 2535 511 2551 545
rect -2597 452 -2563 468
rect -2597 -540 -2563 -524
rect -2339 452 -2305 468
rect -2339 -540 -2305 -524
rect -2081 452 -2047 468
rect -2081 -540 -2047 -524
rect -1823 452 -1789 468
rect -1823 -540 -1789 -524
rect -1565 452 -1531 468
rect -1565 -540 -1531 -524
rect -1307 452 -1273 468
rect -1307 -540 -1273 -524
rect -1049 452 -1015 468
rect -1049 -540 -1015 -524
rect -791 452 -757 468
rect -791 -540 -757 -524
rect -533 452 -499 468
rect -533 -540 -499 -524
rect -275 452 -241 468
rect -275 -540 -241 -524
rect -17 452 17 468
rect -17 -540 17 -524
rect 241 452 275 468
rect 241 -540 275 -524
rect 499 452 533 468
rect 499 -540 533 -524
rect 757 452 791 468
rect 757 -540 791 -524
rect 1015 452 1049 468
rect 1015 -540 1049 -524
rect 1273 452 1307 468
rect 1273 -540 1307 -524
rect 1531 452 1565 468
rect 1531 -540 1565 -524
rect 1789 452 1823 468
rect 1789 -540 1823 -524
rect 2047 452 2081 468
rect 2047 -540 2081 -524
rect 2305 452 2339 468
rect 2305 -540 2339 -524
rect 2563 452 2597 468
rect 2563 -540 2597 -524
rect -2711 -648 -2677 -551
rect 2677 -648 2711 -551
<< viali >>
rect -2493 511 -2409 545
rect -2235 511 -2151 545
rect -1977 511 -1893 545
rect -1719 511 -1635 545
rect -1461 511 -1377 545
rect -1203 511 -1119 545
rect -945 511 -861 545
rect -687 511 -603 545
rect -429 511 -345 545
rect -171 511 -87 545
rect 87 511 171 545
rect 345 511 429 545
rect 603 511 687 545
rect 861 511 945 545
rect 1119 511 1203 545
rect 1377 511 1461 545
rect 1635 511 1719 545
rect 1893 511 1977 545
rect 2151 511 2235 545
rect 2409 511 2493 545
rect -2711 -491 -2677 491
rect -2597 -524 -2563 452
rect -2339 -524 -2305 452
rect -2081 -524 -2047 452
rect -1823 -524 -1789 452
rect -1565 -524 -1531 452
rect -1307 -524 -1273 452
rect -1049 -524 -1015 452
rect -791 -524 -757 452
rect -533 -524 -499 452
rect -275 -524 -241 452
rect -17 -524 17 452
rect 241 -524 275 452
rect 499 -524 533 452
rect 757 -524 791 452
rect 1015 -524 1049 452
rect 1273 -524 1307 452
rect 1531 -524 1565 452
rect 1789 -524 1823 452
rect 2047 -524 2081 452
rect 2305 -524 2339 452
rect 2563 -524 2597 452
rect 2677 -491 2711 491
rect -2677 -648 -2615 -614
rect -2615 -648 2615 -614
rect 2615 -648 2677 -614
<< metal1 >>
rect -2505 545 -2397 551
rect -2505 511 -2493 545
rect -2409 511 -2397 545
rect -2505 505 -2397 511
rect -2247 545 -2139 551
rect -2247 511 -2235 545
rect -2151 511 -2139 545
rect -2247 505 -2139 511
rect -1989 545 -1881 551
rect -1989 511 -1977 545
rect -1893 511 -1881 545
rect -1989 505 -1881 511
rect -1731 545 -1623 551
rect -1731 511 -1719 545
rect -1635 511 -1623 545
rect -1731 505 -1623 511
rect -1473 545 -1365 551
rect -1473 511 -1461 545
rect -1377 511 -1365 545
rect -1473 505 -1365 511
rect -1215 545 -1107 551
rect -1215 511 -1203 545
rect -1119 511 -1107 545
rect -1215 505 -1107 511
rect -957 545 -849 551
rect -957 511 -945 545
rect -861 511 -849 545
rect -957 505 -849 511
rect -699 545 -591 551
rect -699 511 -687 545
rect -603 511 -591 545
rect -699 505 -591 511
rect -441 545 -333 551
rect -441 511 -429 545
rect -345 511 -333 545
rect -441 505 -333 511
rect -183 545 -75 551
rect -183 511 -171 545
rect -87 511 -75 545
rect -183 505 -75 511
rect 75 545 183 551
rect 75 511 87 545
rect 171 511 183 545
rect 75 505 183 511
rect 333 545 441 551
rect 333 511 345 545
rect 429 511 441 545
rect 333 505 441 511
rect 591 545 699 551
rect 591 511 603 545
rect 687 511 699 545
rect 591 505 699 511
rect 849 545 957 551
rect 849 511 861 545
rect 945 511 957 545
rect 849 505 957 511
rect 1107 545 1215 551
rect 1107 511 1119 545
rect 1203 511 1215 545
rect 1107 505 1215 511
rect 1365 545 1473 551
rect 1365 511 1377 545
rect 1461 511 1473 545
rect 1365 505 1473 511
rect 1623 545 1731 551
rect 1623 511 1635 545
rect 1719 511 1731 545
rect 1623 505 1731 511
rect 1881 545 1989 551
rect 1881 511 1893 545
rect 1977 511 1989 545
rect 1881 505 1989 511
rect 2139 545 2247 551
rect 2139 511 2151 545
rect 2235 511 2247 545
rect 2139 505 2247 511
rect 2397 545 2505 551
rect 2397 511 2409 545
rect 2493 511 2505 545
rect 2397 505 2505 511
rect -2717 491 -2671 503
rect -2717 -491 -2711 491
rect -2677 -491 -2671 491
rect 2671 491 2717 503
rect -2717 -503 -2671 -491
rect -2603 452 -2557 464
rect -2603 -524 -2597 452
rect -2563 -524 -2557 452
rect -2603 -536 -2557 -524
rect -2345 452 -2299 464
rect -2345 -524 -2339 452
rect -2305 -524 -2299 452
rect -2345 -536 -2299 -524
rect -2087 452 -2041 464
rect -2087 -524 -2081 452
rect -2047 -524 -2041 452
rect -2087 -536 -2041 -524
rect -1829 452 -1783 464
rect -1829 -524 -1823 452
rect -1789 -524 -1783 452
rect -1829 -536 -1783 -524
rect -1571 452 -1525 464
rect -1571 -524 -1565 452
rect -1531 -524 -1525 452
rect -1571 -536 -1525 -524
rect -1313 452 -1267 464
rect -1313 -524 -1307 452
rect -1273 -524 -1267 452
rect -1313 -536 -1267 -524
rect -1055 452 -1009 464
rect -1055 -524 -1049 452
rect -1015 -524 -1009 452
rect -1055 -536 -1009 -524
rect -797 452 -751 464
rect -797 -524 -791 452
rect -757 -524 -751 452
rect -797 -536 -751 -524
rect -539 452 -493 464
rect -539 -524 -533 452
rect -499 -524 -493 452
rect -539 -536 -493 -524
rect -281 452 -235 464
rect -281 -524 -275 452
rect -241 -524 -235 452
rect -281 -536 -235 -524
rect -23 452 23 464
rect -23 -524 -17 452
rect 17 -524 23 452
rect -23 -536 23 -524
rect 235 452 281 464
rect 235 -524 241 452
rect 275 -524 281 452
rect 235 -536 281 -524
rect 493 452 539 464
rect 493 -524 499 452
rect 533 -524 539 452
rect 493 -536 539 -524
rect 751 452 797 464
rect 751 -524 757 452
rect 791 -524 797 452
rect 751 -536 797 -524
rect 1009 452 1055 464
rect 1009 -524 1015 452
rect 1049 -524 1055 452
rect 1009 -536 1055 -524
rect 1267 452 1313 464
rect 1267 -524 1273 452
rect 1307 -524 1313 452
rect 1267 -536 1313 -524
rect 1525 452 1571 464
rect 1525 -524 1531 452
rect 1565 -524 1571 452
rect 1525 -536 1571 -524
rect 1783 452 1829 464
rect 1783 -524 1789 452
rect 1823 -524 1829 452
rect 1783 -536 1829 -524
rect 2041 452 2087 464
rect 2041 -524 2047 452
rect 2081 -524 2087 452
rect 2041 -536 2087 -524
rect 2299 452 2345 464
rect 2299 -524 2305 452
rect 2339 -524 2345 452
rect 2299 -536 2345 -524
rect 2557 452 2603 464
rect 2557 -524 2563 452
rect 2597 -524 2603 452
rect 2671 -491 2677 491
rect 2711 -491 2717 491
rect 2671 -503 2717 -491
rect 2557 -536 2603 -524
rect -2689 -614 2689 -608
rect -2689 -648 -2677 -614
rect 2677 -648 2689 -614
rect -2689 -654 2689 -648
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -2694 -631 2694 631
string parameters w 5 l 1 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 100 viagr 80 viagl 80 viagt 0
string library sky130
<< end >>
