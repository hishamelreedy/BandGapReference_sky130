magic
tech sky130A
magscale 1 2
timestamp 1634671827
<< nwell >>
rect -4180 326 3034 2473
rect -4180 262 198 326
rect 210 262 3034 326
rect -4180 -2174 3034 262
<< metal1 >>
rect -1946 1524 -1882 1806
rect -1458 1614 -1394 1796
rect -1458 1552 -1268 1614
rect 344 1610 386 1614
rect 458 1610 522 1794
rect 932 1638 996 1798
rect 334 1552 530 1610
rect 672 1558 996 1638
rect -2056 1516 -1858 1524
rect -1794 1516 -1746 1534
rect -2056 1504 -1736 1516
rect -1458 1512 -1394 1552
rect -2060 1478 -1736 1504
rect -2060 1406 -2008 1478
rect -1950 1458 -1736 1478
rect -1594 1484 -1394 1512
rect -1594 1466 -1396 1484
rect -1794 1366 -1746 1458
rect -1588 1396 -1526 1466
rect -1312 1376 -1268 1552
rect -358 1528 -164 1530
rect -1002 1466 148 1528
rect -1794 1338 -1550 1366
rect -842 1356 -796 1374
rect -614 1356 -548 1424
rect -240 1366 -192 1378
rect -1786 1316 -1550 1338
rect -2050 934 -2016 1256
rect -1488 1048 -1386 1056
rect -1488 988 -1464 1048
rect -1406 988 -1386 1048
rect -1488 968 -1386 988
rect -1970 934 -1756 952
rect -2056 928 -1756 934
rect -2056 898 -1750 928
rect -2052 820 -2016 898
rect -1970 894 -1750 898
rect -1808 794 -1750 894
rect -1492 874 -1370 968
rect -1808 756 -1799 794
rect -1790 776 -1562 794
rect -1106 786 -1060 1354
rect -842 1306 -548 1356
rect -328 1314 -100 1366
rect 344 1332 386 1552
rect 458 1482 522 1552
rect 688 1356 756 1558
rect 932 1486 996 1558
rect 1066 1504 1104 1522
rect 1000 1476 1104 1504
rect 1066 1398 1104 1476
rect -312 1312 -288 1314
rect -244 1312 -100 1314
rect -970 1160 -918 1164
rect -984 1048 -912 1160
rect -984 988 -974 1048
rect -916 988 -912 1048
rect -984 972 -912 988
rect -992 888 -906 972
rect -1790 742 -1558 776
rect -1786 724 -1558 742
rect -1298 740 -1060 786
rect -842 794 -796 1306
rect -614 794 -548 1306
rect -470 1072 -418 1170
rect -468 990 -418 1072
rect -472 890 -412 990
rect -842 768 -548 794
rect -240 782 -192 1312
rect 614 1302 826 1356
rect 688 1300 756 1302
rect 10 1072 62 1170
rect 930 1076 982 1174
rect 10 954 60 1072
rect 930 1032 980 1076
rect 1066 1032 1106 1236
rect 802 980 1106 1032
rect 802 970 988 980
rect 422 954 560 966
rect -86 894 560 954
rect -86 882 472 894
rect 526 882 560 894
rect 802 836 850 970
rect 930 906 980 970
rect 1066 832 1106 980
rect -344 780 -192 782
rect -842 760 -566 768
rect -836 744 -566 760
rect -1298 736 -1062 740
rect -2050 418 -2016 712
rect -1930 418 -1880 584
rect -2050 408 -1740 418
rect -2050 368 -1736 408
rect -1446 372 -1398 576
rect -2054 360 -1736 368
rect -2054 356 -1740 360
rect -2054 352 -2016 356
rect -2054 304 -2020 352
rect -1798 292 -1740 356
rect -1798 260 -1738 292
rect -1798 250 -1786 260
rect -1754 250 -1738 260
rect -1802 206 -1538 250
rect -2052 -12 -2018 168
rect -1918 -12 -1870 54
rect -2052 -22 -1844 -12
rect -2052 -74 -1726 -22
rect -2052 -192 -2018 -74
rect -1926 -102 -1726 -74
rect -1440 -100 -1392 52
rect -1320 28 -1274 176
rect -1320 26 -1242 28
rect -1320 -50 -1314 26
rect -1250 -50 -1242 26
rect -1320 -60 -1242 -50
rect -1320 -64 -1274 -60
rect -1918 -150 -1870 -102
rect -2050 -226 -2020 -192
rect -1780 -282 -1732 -102
rect -1444 -158 -1386 -100
rect -1208 -130 -1172 736
rect -964 384 -916 588
rect -836 252 -798 744
rect -738 370 -656 378
rect -738 296 -728 370
rect -748 280 -728 296
rect -668 280 -656 370
rect -748 252 -656 280
rect -600 252 -566 744
rect -344 730 -90 780
rect 142 732 400 782
rect 596 774 752 778
rect -344 726 -192 730
rect -240 714 -192 726
rect -464 398 -416 582
rect -464 378 -290 398
rect -416 358 -290 378
rect -344 276 -294 358
rect -836 202 -566 252
rect -1090 40 -1048 166
rect -836 138 -798 202
rect -748 196 -656 202
rect -1140 18 -1042 40
rect -1140 -58 -1118 18
rect -1054 -58 -1042 18
rect -1140 -76 -1042 -58
rect -962 -96 -914 50
rect -970 -154 -912 -96
rect -748 -146 -660 196
rect -600 174 -566 202
rect -480 -142 -432 62
rect -342 58 -296 184
rect -352 54 -284 58
rect -354 44 -278 54
rect -290 -32 -278 44
rect -354 -68 -278 -32
rect -1208 -282 -1172 -178
rect -752 -230 -660 -146
rect -752 -246 -590 -230
rect -1800 -346 -1526 -282
rect -1304 -332 -1068 -282
rect -824 -300 -590 -246
rect -824 -304 -668 -300
rect -2054 -590 -2014 -388
rect -1780 -398 -1732 -346
rect -1208 -410 -1142 -332
rect -1920 -590 -1872 -488
rect -2070 -622 -1860 -590
rect -2054 -792 -2014 -622
rect -1920 -686 -1872 -622
rect -1560 -676 -1516 -672
rect -1412 -676 -1254 -666
rect -1692 -686 -1638 -680
rect -1920 -692 -1638 -686
rect -1890 -716 -1638 -692
rect -1692 -816 -1638 -716
rect -1560 -718 -1254 -676
rect -1560 -800 -1516 -718
rect -1298 -790 -1256 -718
rect -1782 -866 -1546 -816
rect -1198 -840 -1142 -410
rect -980 -508 -918 -482
rect -980 -616 -914 -508
rect -968 -706 -914 -616
rect -752 -806 -668 -304
rect -566 -542 -472 -534
rect -566 -602 -560 -542
rect -502 -544 -472 -542
rect -372 -544 -318 -268
rect -502 -592 -318 -544
rect -502 -602 -320 -592
rect -566 -606 -320 -602
rect -566 -614 -472 -606
rect -486 -706 -440 -692
rect -1206 -920 -1052 -840
rect -832 -872 -582 -806
rect -236 -808 -192 714
rect 14 388 62 592
rect 142 264 194 732
rect 596 728 758 774
rect 224 482 286 486
rect 224 478 294 482
rect 224 418 230 478
rect 288 418 294 478
rect 224 362 294 418
rect 474 374 522 578
rect 226 264 294 362
rect 142 262 198 264
rect 226 262 378 264
rect 140 214 378 262
rect 232 210 292 214
rect -122 46 -70 162
rect -144 38 -70 46
rect -144 30 -56 38
rect -144 -46 -132 30
rect -68 -46 -56 30
rect -144 -54 -56 -46
rect -144 -66 -78 -54
rect 14 -130 62 64
rect 232 -30 282 210
rect 594 72 642 146
rect 228 -130 282 -30
rect 464 -130 512 54
rect 592 30 672 72
rect 592 -46 600 30
rect 664 -46 672 30
rect 592 -66 672 -46
rect 228 -178 278 -130
rect 228 -226 282 -178
rect -256 -812 -176 -808
rect -148 -812 -88 -234
rect 232 -258 282 -226
rect 716 -242 758 728
rect 932 522 980 588
rect 1072 522 1112 688
rect 806 502 850 522
rect 932 502 1116 522
rect 796 470 1116 502
rect 796 456 992 470
rect 806 250 850 456
rect 932 384 980 456
rect 1072 284 1112 470
rect 938 -32 986 56
rect 1068 -32 1108 162
rect 938 -84 1116 -32
rect 938 -118 986 -84
rect 812 -128 986 -118
rect 142 -308 378 -258
rect 592 -366 758 -242
rect 806 -148 986 -128
rect 806 -170 978 -148
rect 806 -280 848 -170
rect 1068 -242 1108 -84
rect 6 -670 54 -498
rect 210 -524 322 -514
rect 210 -600 234 -524
rect 298 -544 322 -524
rect 604 -544 636 -366
rect 298 -576 636 -544
rect 940 -552 988 -478
rect 1078 -552 1118 -366
rect 298 -600 634 -576
rect 210 -622 322 -600
rect 940 -604 1118 -552
rect 940 -654 988 -604
rect 330 -678 548 -660
rect 330 -706 654 -678
rect 818 -682 988 -654
rect 818 -702 960 -682
rect 330 -714 548 -706
rect 338 -790 396 -714
rect 614 -764 654 -706
rect 820 -748 860 -702
rect 1078 -770 1118 -604
rect -348 -880 -88 -812
rect -348 -896 -110 -880
rect -252 -898 -110 -896
rect -1202 -1406 -1146 -920
rect -236 -936 -192 -898
rect 168 -900 378 -836
rect 610 -862 846 -812
rect -994 -1044 -424 -1000
rect -236 -1398 -194 -936
rect 214 -1062 300 -1038
rect 214 -1138 230 -1062
rect 294 -1130 300 -1062
rect 294 -1138 302 -1130
rect 214 -1360 302 -1138
rect 216 -1398 302 -1360
rect -790 -1406 -580 -1402
rect -260 -1406 302 -1398
rect -1202 -1462 302 -1406
rect -1202 -1464 -194 -1462
rect -790 -1472 -580 -1464
<< via1 >>
rect -1464 988 -1406 1048
rect -974 988 -916 1048
rect -1314 -50 -1250 26
rect -728 280 -668 370
rect -1118 -58 -1054 18
rect -354 -32 -290 44
rect -560 -602 -502 -542
rect 230 418 288 478
rect -132 -46 -68 30
rect 600 -46 664 30
rect 234 -600 298 -524
rect 230 -1138 294 -1062
<< metal2 >>
rect -2396 1808 1483 1852
rect -2396 1724 -746 1808
rect -664 1724 220 1808
rect 302 1724 1483 1808
rect -2396 1710 1483 1724
rect -940 1056 -912 1058
rect -1490 1048 -912 1056
rect -1490 988 -1464 1048
rect -1406 988 -974 1048
rect -916 988 -912 1048
rect -1490 976 -912 988
rect -940 974 -912 976
rect 208 628 302 644
rect -746 564 -658 576
rect -746 466 -728 564
rect -662 466 -658 564
rect 208 530 224 628
rect 290 530 302 628
rect 208 516 302 530
rect -746 432 -658 466
rect 228 478 294 516
rect -746 424 -660 432
rect -740 370 -660 424
rect 228 418 230 478
rect 288 418 294 478
rect 228 410 294 418
rect 228 408 290 410
rect -740 280 -728 370
rect -668 280 -660 370
rect -740 270 -660 280
rect -320 58 -278 60
rect -352 54 -278 58
rect -352 52 -250 54
rect -356 44 -250 52
rect -1322 26 -1244 38
rect -1322 -50 -1314 26
rect -1250 -50 -1244 26
rect -1322 -108 -1244 -50
rect -1140 34 -1042 40
rect -1140 18 -1038 34
rect -1140 -58 -1118 18
rect -1054 -58 -1038 18
rect -1140 -68 -1038 -58
rect -356 -32 -354 44
rect -290 -32 -250 44
rect -1140 -76 -1042 -68
rect -356 -72 -250 -32
rect -178 30 -56 54
rect -178 -46 -132 30
rect -68 -46 -56 30
rect -178 -54 -56 -46
rect 578 30 670 56
rect 578 -46 600 30
rect 664 -46 670 30
rect -1310 -314 -1266 -108
rect -1136 -166 -1088 -76
rect -1310 -1152 -1262 -314
rect -1134 -1114 -1090 -166
rect -746 -542 -490 -532
rect -746 -602 -560 -542
rect -502 -602 -490 -542
rect -746 -618 -490 -602
rect -746 -1082 -662 -618
rect -1306 -1278 -1262 -1152
rect -1310 -1444 -1262 -1278
rect -1140 -1182 -1090 -1114
rect -1140 -1336 -1094 -1182
rect -750 -1232 -660 -1082
rect -352 -1104 -308 -72
rect -178 -76 -62 -54
rect 578 -72 670 -46
rect -178 -78 -90 -76
rect -134 -1032 -90 -78
rect -362 -1182 -308 -1104
rect -140 -1180 -90 -1032
rect 220 -524 304 -520
rect 220 -600 234 -524
rect 298 -600 304 -524
rect 220 -1062 304 -600
rect 220 -1138 230 -1062
rect 294 -1138 304 -1062
rect 220 -1156 304 -1138
rect -1310 -1886 -1264 -1444
rect -1146 -1722 -1094 -1336
rect -362 -1412 -316 -1182
rect -368 -1712 -316 -1412
rect -140 -1388 -94 -1180
rect 578 -1356 680 -72
rect -140 -1640 -90 -1388
rect 578 -1496 684 -1356
rect -1146 -1944 -1100 -1722
rect -368 -2020 -322 -1712
rect -136 -1996 -90 -1640
rect 586 -1948 684 -1496
<< via2 >>
rect -746 1724 -664 1808
rect 220 1724 302 1808
rect -728 466 -662 564
rect 224 530 290 628
<< metal3 >>
rect -758 1808 -658 1816
rect -758 1724 -746 1808
rect -664 1724 -658 1808
rect -758 1712 -658 1724
rect -746 598 -658 1712
rect 210 1808 310 1814
rect 210 1724 220 1808
rect 302 1724 310 1808
rect 210 1708 310 1724
rect 224 640 300 1708
rect 216 638 300 640
rect 216 628 304 638
rect 216 626 224 628
rect -748 564 -654 598
rect -748 466 -728 564
rect -662 466 -654 564
rect 214 530 224 626
rect 290 530 304 628
rect 214 524 304 530
rect 214 520 296 524
rect -748 454 -654 466
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_7
timestamp 1634549143
transform 1 0 -1908 0 1 -859
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_12
timestamp 1634505583
transform 1 0 -943 0 1 -861
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_13
timestamp 1634549143
transform 1 0 -1408 0 1 -861
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_13
timestamp 1634505583
transform 1 0 -472 0 1 -857
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_14
timestamp 1634505583
transform 1 0 16 0 1 -856
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_12
timestamp 1634549143
transform 1 0 501 0 1 -857
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_11
timestamp 1634549143
transform 1 0 967 0 1 -841
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_6
timestamp 1634549143
transform 1 0 -1901 0 1 -320
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_10
timestamp 1634505583
transform 1 0 -940 0 1 -322
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_11
timestamp 1634505583
transform 1 0 -1413 0 1 -320
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M12  sky130_fd_pr__pfet_01v8_lvt_M12_0
timestamp 1634505583
transform 1 0 -472 0 1 -314
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_9
timestamp 1634505583
transform 1 0 34 0 1 -313
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_8
timestamp 1634505583
transform 1 0 493 0 1 -316
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_10
timestamp 1634549143
transform 1 0 957 0 1 -318
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_5
timestamp 1634549143
transform 1 0 -1905 0 1 219
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M11  sky130_fd_pr__pfet_01v8_lvt_M11_0
timestamp 1634505583
transform 1 0 -1426 0 1 221
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M10  sky130_fd_pr__pfet_01v8_lvt_M10_0
timestamp 1634505583
transform 1 0 -940 0 1 223
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M8  sky130_fd_pr__pfet_01v8_lvt_M8_0
timestamp 1634505583
transform 1 0 -449 0 1 218
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M13  sky130_fd_pr__pfet_01v8_lvt_M13_0
timestamp 1634505583
transform 1 0 34 0 1 227
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M16  sky130_fd_pr__pfet_01v8_lvt_M16_0
timestamp 1634505583
transform 1 0 491 0 1 214
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_8
timestamp 1634549143
transform 1 0 957 0 1 218
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_4
timestamp 1634549143
transform 1 0 -1905 0 1 747
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_3
timestamp 1634505583
transform 1 0 -1428 0 1 740
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_4
timestamp 1634505583
transform 1 0 -946 0 1 744
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_5
timestamp 1634505583
transform 1 0 -447 0 1 742
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_6
timestamp 1634505583
transform 1 0 37 0 1 744
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_7
timestamp 1634505583
transform 1 0 496 0 1 744
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_9
timestamp 1634549143
transform 1 0 957 0 1 751
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_3
timestamp 1634549143
transform 1 0 -1905 0 1 1324
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_2
timestamp 1634549143
transform 1 0 -1424 0 1 1321
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_0
timestamp 1634505583
transform -1 0 -947 0 1 1322
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_1
timestamp 1634505583
transform 1 0 -443 0 1 1324
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_M9  sky130_fd_pr__pfet_01v8_lvt_M9_2
timestamp 1634505583
transform 1 0 32 0 1 1322
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_0
timestamp 1634549143
transform 1 0 494 0 1 1321
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_lvt_MD  sky130_fd_pr__pfet_01v8_lvt_MD_1
timestamp 1634549143
transform 1 0 957 0 1 1326
box -194 -200 194 200
<< labels >>
flabel metal2 -2396 1710 1483 1852 0 FreeSans 1600 0 0 0 VDD
flabel metal2 586 -1948 684 -1356 0 FreeSans 800 0 0 0 M16D
flabel metal2 -136 -1996 -90 -1388 0 FreeSans 800 0 0 0 M13D
flabel metal2 -368 -2020 -322 -1412 0 FreeSans 800 0 0 0 M8D
flabel metal2 -1146 -1944 -1100 -1336 0 FreeSans 800 0 0 0 M10D
flabel metal2 -1310 -1886 -1264 -1278 0 FreeSans 800 0 0 0 M11D
flabel metal2 -750 -1232 -660 -1082 0 FreeSans 480 0 0 0 M12D
<< end >>
