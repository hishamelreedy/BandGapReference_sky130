magic
tech sky130A
magscale 1 2
timestamp 1629311173
<< checkpaint >>
rect -1260 -1260 5758 3598
<< poly >>
rect 0 2322 4498 2338
rect 0 2288 34 2322
rect 68 2288 102 2322
rect 136 2288 170 2322
rect 204 2288 238 2322
rect 272 2288 306 2322
rect 340 2288 374 2322
rect 408 2288 442 2322
rect 476 2288 510 2322
rect 544 2288 578 2322
rect 612 2288 646 2322
rect 680 2288 714 2322
rect 748 2288 782 2322
rect 816 2288 850 2322
rect 884 2288 918 2322
rect 952 2288 986 2322
rect 1020 2288 1054 2322
rect 1088 2288 1122 2322
rect 1156 2288 1190 2322
rect 1224 2288 1258 2322
rect 1292 2288 1326 2322
rect 1360 2288 1394 2322
rect 1428 2288 1462 2322
rect 1496 2288 1530 2322
rect 1564 2288 1598 2322
rect 1632 2288 1666 2322
rect 1700 2288 1734 2322
rect 1768 2288 1802 2322
rect 1836 2288 1870 2322
rect 1904 2288 1938 2322
rect 1972 2288 2006 2322
rect 2040 2288 2074 2322
rect 2108 2288 2142 2322
rect 2176 2288 2210 2322
rect 2244 2288 2278 2322
rect 2312 2288 2346 2322
rect 2380 2288 2414 2322
rect 2448 2288 2482 2322
rect 2516 2288 2550 2322
rect 2584 2288 2618 2322
rect 2652 2288 2686 2322
rect 2720 2288 2754 2322
rect 2788 2288 2822 2322
rect 2856 2288 2890 2322
rect 2924 2288 2958 2322
rect 2992 2288 3026 2322
rect 3060 2288 3094 2322
rect 3128 2288 3162 2322
rect 3196 2288 3230 2322
rect 3264 2288 3298 2322
rect 3332 2288 3366 2322
rect 3400 2288 3434 2322
rect 3468 2288 3502 2322
rect 3536 2288 3570 2322
rect 3604 2288 3638 2322
rect 3672 2288 3706 2322
rect 3740 2288 3774 2322
rect 3808 2288 3842 2322
rect 3876 2288 3910 2322
rect 3944 2288 3978 2322
rect 4012 2288 4046 2322
rect 4080 2288 4114 2322
rect 4148 2288 4182 2322
rect 4216 2288 4250 2322
rect 4284 2288 4318 2322
rect 4352 2288 4386 2322
rect 4420 2288 4498 2322
rect 0 2272 4498 2288
rect 0 108 30 2272
rect 72 66 102 2230
rect 144 108 174 2272
rect 216 66 246 2230
rect 288 108 318 2272
rect 360 66 390 2230
rect 432 108 462 2272
rect 504 66 534 2230
rect 576 108 606 2272
rect 648 66 678 2230
rect 720 108 750 2272
rect 792 66 822 2230
rect 864 108 894 2272
rect 936 66 966 2230
rect 1008 108 1038 2272
rect 1080 66 1110 2230
rect 1152 108 1182 2272
rect 1224 66 1254 2230
rect 1296 108 1326 2272
rect 1368 66 1398 2230
rect 1440 108 1470 2272
rect 1512 66 1542 2230
rect 1584 108 1614 2272
rect 1656 66 1686 2230
rect 1728 108 1758 2272
rect 1800 66 1830 2230
rect 1872 108 1902 2272
rect 1944 66 1974 2230
rect 2016 108 2046 2272
rect 2088 66 2118 2230
rect 2160 108 2190 2272
rect 2232 66 2262 2230
rect 2304 108 2334 2272
rect 2376 66 2406 2230
rect 2448 108 2478 2272
rect 2520 66 2550 2230
rect 2592 108 2622 2272
rect 2664 66 2694 2230
rect 2736 108 2766 2272
rect 2808 66 2838 2230
rect 2880 108 2910 2272
rect 2952 66 2982 2230
rect 3024 108 3054 2272
rect 3096 66 3126 2230
rect 3168 108 3198 2272
rect 3240 66 3270 2230
rect 3312 108 3342 2272
rect 3384 66 3414 2230
rect 3456 108 3486 2272
rect 3528 66 3558 2230
rect 3600 108 3630 2272
rect 3672 66 3702 2230
rect 3744 108 3774 2272
rect 3816 66 3846 2230
rect 3888 108 3918 2272
rect 3960 66 3990 2230
rect 4032 108 4062 2272
rect 4104 66 4134 2230
rect 4176 108 4206 2272
rect 4248 66 4278 2230
rect 4320 108 4350 2272
rect 4392 66 4422 2230
rect 4464 108 4498 2272
rect 0 50 4498 66
rect 0 16 34 50
rect 68 16 102 50
rect 136 16 170 50
rect 204 16 238 50
rect 272 16 306 50
rect 340 16 374 50
rect 408 16 442 50
rect 476 16 510 50
rect 544 16 578 50
rect 612 16 646 50
rect 680 16 714 50
rect 748 16 782 50
rect 816 16 850 50
rect 884 16 918 50
rect 952 16 986 50
rect 1020 16 1054 50
rect 1088 16 1122 50
rect 1156 16 1190 50
rect 1224 16 1258 50
rect 1292 16 1326 50
rect 1360 16 1394 50
rect 1428 16 1462 50
rect 1496 16 1530 50
rect 1564 16 1598 50
rect 1632 16 1666 50
rect 1700 16 1734 50
rect 1768 16 1802 50
rect 1836 16 1870 50
rect 1904 16 1938 50
rect 1972 16 2006 50
rect 2040 16 2074 50
rect 2108 16 2142 50
rect 2176 16 2210 50
rect 2244 16 2278 50
rect 2312 16 2346 50
rect 2380 16 2414 50
rect 2448 16 2482 50
rect 2516 16 2550 50
rect 2584 16 2618 50
rect 2652 16 2686 50
rect 2720 16 2754 50
rect 2788 16 2822 50
rect 2856 16 2890 50
rect 2924 16 2958 50
rect 2992 16 3026 50
rect 3060 16 3094 50
rect 3128 16 3162 50
rect 3196 16 3230 50
rect 3264 16 3298 50
rect 3332 16 3366 50
rect 3400 16 3434 50
rect 3468 16 3502 50
rect 3536 16 3570 50
rect 3604 16 3638 50
rect 3672 16 3706 50
rect 3740 16 3774 50
rect 3808 16 3842 50
rect 3876 16 3910 50
rect 3944 16 3978 50
rect 4012 16 4046 50
rect 4080 16 4114 50
rect 4148 16 4182 50
rect 4216 16 4250 50
rect 4284 16 4318 50
rect 4352 16 4386 50
rect 4420 16 4498 50
rect 0 0 4498 16
<< polycont >>
rect 34 2288 68 2322
rect 102 2288 136 2322
rect 170 2288 204 2322
rect 238 2288 272 2322
rect 306 2288 340 2322
rect 374 2288 408 2322
rect 442 2288 476 2322
rect 510 2288 544 2322
rect 578 2288 612 2322
rect 646 2288 680 2322
rect 714 2288 748 2322
rect 782 2288 816 2322
rect 850 2288 884 2322
rect 918 2288 952 2322
rect 986 2288 1020 2322
rect 1054 2288 1088 2322
rect 1122 2288 1156 2322
rect 1190 2288 1224 2322
rect 1258 2288 1292 2322
rect 1326 2288 1360 2322
rect 1394 2288 1428 2322
rect 1462 2288 1496 2322
rect 1530 2288 1564 2322
rect 1598 2288 1632 2322
rect 1666 2288 1700 2322
rect 1734 2288 1768 2322
rect 1802 2288 1836 2322
rect 1870 2288 1904 2322
rect 1938 2288 1972 2322
rect 2006 2288 2040 2322
rect 2074 2288 2108 2322
rect 2142 2288 2176 2322
rect 2210 2288 2244 2322
rect 2278 2288 2312 2322
rect 2346 2288 2380 2322
rect 2414 2288 2448 2322
rect 2482 2288 2516 2322
rect 2550 2288 2584 2322
rect 2618 2288 2652 2322
rect 2686 2288 2720 2322
rect 2754 2288 2788 2322
rect 2822 2288 2856 2322
rect 2890 2288 2924 2322
rect 2958 2288 2992 2322
rect 3026 2288 3060 2322
rect 3094 2288 3128 2322
rect 3162 2288 3196 2322
rect 3230 2288 3264 2322
rect 3298 2288 3332 2322
rect 3366 2288 3400 2322
rect 3434 2288 3468 2322
rect 3502 2288 3536 2322
rect 3570 2288 3604 2322
rect 3638 2288 3672 2322
rect 3706 2288 3740 2322
rect 3774 2288 3808 2322
rect 3842 2288 3876 2322
rect 3910 2288 3944 2322
rect 3978 2288 4012 2322
rect 4046 2288 4080 2322
rect 4114 2288 4148 2322
rect 4182 2288 4216 2322
rect 4250 2288 4284 2322
rect 4318 2288 4352 2322
rect 4386 2288 4420 2322
rect 34 16 68 50
rect 102 16 136 50
rect 170 16 204 50
rect 238 16 272 50
rect 306 16 340 50
rect 374 16 408 50
rect 442 16 476 50
rect 510 16 544 50
rect 578 16 612 50
rect 646 16 680 50
rect 714 16 748 50
rect 782 16 816 50
rect 850 16 884 50
rect 918 16 952 50
rect 986 16 1020 50
rect 1054 16 1088 50
rect 1122 16 1156 50
rect 1190 16 1224 50
rect 1258 16 1292 50
rect 1326 16 1360 50
rect 1394 16 1428 50
rect 1462 16 1496 50
rect 1530 16 1564 50
rect 1598 16 1632 50
rect 1666 16 1700 50
rect 1734 16 1768 50
rect 1802 16 1836 50
rect 1870 16 1904 50
rect 1938 16 1972 50
rect 2006 16 2040 50
rect 2074 16 2108 50
rect 2142 16 2176 50
rect 2210 16 2244 50
rect 2278 16 2312 50
rect 2346 16 2380 50
rect 2414 16 2448 50
rect 2482 16 2516 50
rect 2550 16 2584 50
rect 2618 16 2652 50
rect 2686 16 2720 50
rect 2754 16 2788 50
rect 2822 16 2856 50
rect 2890 16 2924 50
rect 2958 16 2992 50
rect 3026 16 3060 50
rect 3094 16 3128 50
rect 3162 16 3196 50
rect 3230 16 3264 50
rect 3298 16 3332 50
rect 3366 16 3400 50
rect 3434 16 3468 50
rect 3502 16 3536 50
rect 3570 16 3604 50
rect 3638 16 3672 50
rect 3706 16 3740 50
rect 3774 16 3808 50
rect 3842 16 3876 50
rect 3910 16 3944 50
rect 3978 16 4012 50
rect 4046 16 4080 50
rect 4114 16 4148 50
rect 4182 16 4216 50
rect 4250 16 4284 50
rect 4318 16 4352 50
rect 4386 16 4420 50
<< locali >>
rect 0 2322 4498 2338
rect 0 2288 34 2322
rect 72 2288 102 2322
rect 144 2288 170 2322
rect 216 2288 238 2322
rect 288 2288 306 2322
rect 360 2288 374 2322
rect 432 2288 442 2322
rect 504 2288 510 2322
rect 576 2288 578 2322
rect 612 2288 614 2322
rect 680 2288 686 2322
rect 748 2288 758 2322
rect 816 2288 830 2322
rect 884 2288 902 2322
rect 952 2288 974 2322
rect 1020 2288 1046 2322
rect 1088 2288 1118 2322
rect 1156 2288 1190 2322
rect 1224 2288 1258 2322
rect 1296 2288 1326 2322
rect 1368 2288 1394 2322
rect 1440 2288 1462 2322
rect 1512 2288 1530 2322
rect 1584 2288 1598 2322
rect 1656 2288 1666 2322
rect 1728 2288 1734 2322
rect 1800 2288 1802 2322
rect 1836 2288 1838 2322
rect 1904 2288 1910 2322
rect 1972 2288 1982 2322
rect 2040 2288 2054 2322
rect 2108 2288 2126 2322
rect 2176 2288 2198 2322
rect 2244 2288 2270 2322
rect 2312 2288 2342 2322
rect 2380 2288 2414 2322
rect 2448 2288 2482 2322
rect 2520 2288 2550 2322
rect 2592 2288 2618 2322
rect 2664 2288 2686 2322
rect 2736 2288 2754 2322
rect 2808 2288 2822 2322
rect 2880 2288 2890 2322
rect 2952 2288 2958 2322
rect 3024 2288 3026 2322
rect 3060 2288 3062 2322
rect 3128 2288 3134 2322
rect 3196 2288 3206 2322
rect 3264 2288 3278 2322
rect 3332 2288 3350 2322
rect 3400 2288 3422 2322
rect 3468 2288 3494 2322
rect 3536 2288 3566 2322
rect 3604 2288 3638 2322
rect 3672 2288 3706 2322
rect 3744 2288 3774 2322
rect 3816 2288 3842 2322
rect 3888 2288 3910 2322
rect 3960 2288 3978 2322
rect 4032 2288 4046 2322
rect 4104 2288 4114 2322
rect 4176 2288 4182 2322
rect 4248 2288 4250 2322
rect 4284 2288 4286 2322
rect 4352 2288 4358 2322
rect 4420 2288 4498 2322
rect 0 2272 4498 2288
rect 0 66 28 2244
rect 56 94 84 2272
rect 112 66 140 2244
rect 168 94 196 2272
rect 224 66 252 2244
rect 280 94 308 2272
rect 336 66 364 2244
rect 392 94 420 2272
rect 448 66 476 2244
rect 504 94 532 2272
rect 560 66 588 2244
rect 616 94 644 2272
rect 672 66 700 2244
rect 728 94 756 2272
rect 784 66 812 2244
rect 840 94 868 2272
rect 896 66 924 2244
rect 952 94 980 2272
rect 1008 66 1036 2244
rect 1064 94 1092 2272
rect 1120 66 1148 2244
rect 1176 94 1204 2272
rect 1232 66 1260 2244
rect 1288 94 1316 2272
rect 1344 66 1372 2244
rect 1400 94 1428 2272
rect 1456 66 1484 2244
rect 1512 94 1540 2272
rect 1568 66 1596 2244
rect 1624 94 1652 2272
rect 1680 66 1708 2244
rect 1736 94 1764 2272
rect 1792 66 1820 2244
rect 1848 94 1876 2272
rect 1904 66 1932 2244
rect 1960 94 1988 2272
rect 2016 66 2044 2244
rect 2072 94 2100 2272
rect 2128 66 2156 2244
rect 2184 94 2212 2272
rect 2240 66 2268 2244
rect 2296 94 2324 2272
rect 2352 66 2380 2244
rect 2408 94 2436 2272
rect 2464 66 2492 2244
rect 2520 94 2548 2272
rect 2576 66 2604 2244
rect 2632 94 2660 2272
rect 2688 66 2716 2244
rect 2744 94 2772 2272
rect 2800 66 2828 2244
rect 2856 94 2884 2272
rect 2912 66 2940 2244
rect 2968 94 2996 2272
rect 3024 66 3052 2244
rect 3080 94 3108 2272
rect 3136 66 3164 2244
rect 3192 94 3220 2272
rect 3248 66 3276 2244
rect 3304 94 3332 2272
rect 3360 66 3388 2244
rect 3416 94 3444 2272
rect 3472 66 3500 2244
rect 3528 94 3556 2272
rect 3584 66 3612 2244
rect 3640 94 3668 2272
rect 3696 66 3724 2244
rect 3752 94 3780 2272
rect 3808 66 3836 2244
rect 3864 94 3892 2272
rect 3920 66 3948 2244
rect 3976 94 4004 2272
rect 4032 66 4060 2244
rect 4088 94 4116 2272
rect 4144 66 4172 2244
rect 4200 94 4228 2272
rect 4256 66 4284 2244
rect 4312 94 4340 2272
rect 4368 66 4396 2244
rect 4424 94 4498 2272
rect 0 50 4498 66
rect 0 16 34 50
rect 72 16 102 50
rect 144 16 170 50
rect 216 16 238 50
rect 288 16 306 50
rect 360 16 374 50
rect 432 16 442 50
rect 504 16 510 50
rect 576 16 578 50
rect 612 16 614 50
rect 680 16 686 50
rect 748 16 758 50
rect 816 16 830 50
rect 884 16 902 50
rect 952 16 974 50
rect 1020 16 1046 50
rect 1088 16 1118 50
rect 1156 16 1190 50
rect 1224 16 1258 50
rect 1296 16 1326 50
rect 1368 16 1394 50
rect 1440 16 1462 50
rect 1512 16 1530 50
rect 1584 16 1598 50
rect 1656 16 1666 50
rect 1728 16 1734 50
rect 1800 16 1802 50
rect 1836 16 1838 50
rect 1904 16 1910 50
rect 1972 16 1982 50
rect 2040 16 2054 50
rect 2108 16 2126 50
rect 2176 16 2198 50
rect 2244 16 2270 50
rect 2312 16 2342 50
rect 2380 16 2414 50
rect 2448 16 2482 50
rect 2520 16 2550 50
rect 2592 16 2618 50
rect 2664 16 2686 50
rect 2736 16 2754 50
rect 2808 16 2822 50
rect 2880 16 2890 50
rect 2952 16 2958 50
rect 3024 16 3026 50
rect 3060 16 3062 50
rect 3128 16 3134 50
rect 3196 16 3206 50
rect 3264 16 3278 50
rect 3332 16 3350 50
rect 3400 16 3422 50
rect 3468 16 3494 50
rect 3536 16 3566 50
rect 3604 16 3638 50
rect 3672 16 3706 50
rect 3744 16 3774 50
rect 3816 16 3842 50
rect 3888 16 3910 50
rect 3960 16 3978 50
rect 4032 16 4046 50
rect 4104 16 4114 50
rect 4176 16 4182 50
rect 4248 16 4250 50
rect 4284 16 4286 50
rect 4352 16 4358 50
rect 4420 16 4498 50
rect 0 0 4498 16
<< viali >>
rect 38 2288 68 2322
rect 68 2288 72 2322
rect 110 2288 136 2322
rect 136 2288 144 2322
rect 182 2288 204 2322
rect 204 2288 216 2322
rect 254 2288 272 2322
rect 272 2288 288 2322
rect 326 2288 340 2322
rect 340 2288 360 2322
rect 398 2288 408 2322
rect 408 2288 432 2322
rect 470 2288 476 2322
rect 476 2288 504 2322
rect 542 2288 544 2322
rect 544 2288 576 2322
rect 614 2288 646 2322
rect 646 2288 648 2322
rect 686 2288 714 2322
rect 714 2288 720 2322
rect 758 2288 782 2322
rect 782 2288 792 2322
rect 830 2288 850 2322
rect 850 2288 864 2322
rect 902 2288 918 2322
rect 918 2288 936 2322
rect 974 2288 986 2322
rect 986 2288 1008 2322
rect 1046 2288 1054 2322
rect 1054 2288 1080 2322
rect 1118 2288 1122 2322
rect 1122 2288 1152 2322
rect 1190 2288 1224 2322
rect 1262 2288 1292 2322
rect 1292 2288 1296 2322
rect 1334 2288 1360 2322
rect 1360 2288 1368 2322
rect 1406 2288 1428 2322
rect 1428 2288 1440 2322
rect 1478 2288 1496 2322
rect 1496 2288 1512 2322
rect 1550 2288 1564 2322
rect 1564 2288 1584 2322
rect 1622 2288 1632 2322
rect 1632 2288 1656 2322
rect 1694 2288 1700 2322
rect 1700 2288 1728 2322
rect 1766 2288 1768 2322
rect 1768 2288 1800 2322
rect 1838 2288 1870 2322
rect 1870 2288 1872 2322
rect 1910 2288 1938 2322
rect 1938 2288 1944 2322
rect 1982 2288 2006 2322
rect 2006 2288 2016 2322
rect 2054 2288 2074 2322
rect 2074 2288 2088 2322
rect 2126 2288 2142 2322
rect 2142 2288 2160 2322
rect 2198 2288 2210 2322
rect 2210 2288 2232 2322
rect 2270 2288 2278 2322
rect 2278 2288 2304 2322
rect 2342 2288 2346 2322
rect 2346 2288 2376 2322
rect 2414 2288 2448 2322
rect 2486 2288 2516 2322
rect 2516 2288 2520 2322
rect 2558 2288 2584 2322
rect 2584 2288 2592 2322
rect 2630 2288 2652 2322
rect 2652 2288 2664 2322
rect 2702 2288 2720 2322
rect 2720 2288 2736 2322
rect 2774 2288 2788 2322
rect 2788 2288 2808 2322
rect 2846 2288 2856 2322
rect 2856 2288 2880 2322
rect 2918 2288 2924 2322
rect 2924 2288 2952 2322
rect 2990 2288 2992 2322
rect 2992 2288 3024 2322
rect 3062 2288 3094 2322
rect 3094 2288 3096 2322
rect 3134 2288 3162 2322
rect 3162 2288 3168 2322
rect 3206 2288 3230 2322
rect 3230 2288 3240 2322
rect 3278 2288 3298 2322
rect 3298 2288 3312 2322
rect 3350 2288 3366 2322
rect 3366 2288 3384 2322
rect 3422 2288 3434 2322
rect 3434 2288 3456 2322
rect 3494 2288 3502 2322
rect 3502 2288 3528 2322
rect 3566 2288 3570 2322
rect 3570 2288 3600 2322
rect 3638 2288 3672 2322
rect 3710 2288 3740 2322
rect 3740 2288 3744 2322
rect 3782 2288 3808 2322
rect 3808 2288 3816 2322
rect 3854 2288 3876 2322
rect 3876 2288 3888 2322
rect 3926 2288 3944 2322
rect 3944 2288 3960 2322
rect 3998 2288 4012 2322
rect 4012 2288 4032 2322
rect 4070 2288 4080 2322
rect 4080 2288 4104 2322
rect 4142 2288 4148 2322
rect 4148 2288 4176 2322
rect 4214 2288 4216 2322
rect 4216 2288 4248 2322
rect 4286 2288 4318 2322
rect 4318 2288 4320 2322
rect 4358 2288 4386 2322
rect 4386 2288 4392 2322
rect 38 16 68 50
rect 68 16 72 50
rect 110 16 136 50
rect 136 16 144 50
rect 182 16 204 50
rect 204 16 216 50
rect 254 16 272 50
rect 272 16 288 50
rect 326 16 340 50
rect 340 16 360 50
rect 398 16 408 50
rect 408 16 432 50
rect 470 16 476 50
rect 476 16 504 50
rect 542 16 544 50
rect 544 16 576 50
rect 614 16 646 50
rect 646 16 648 50
rect 686 16 714 50
rect 714 16 720 50
rect 758 16 782 50
rect 782 16 792 50
rect 830 16 850 50
rect 850 16 864 50
rect 902 16 918 50
rect 918 16 936 50
rect 974 16 986 50
rect 986 16 1008 50
rect 1046 16 1054 50
rect 1054 16 1080 50
rect 1118 16 1122 50
rect 1122 16 1152 50
rect 1190 16 1224 50
rect 1262 16 1292 50
rect 1292 16 1296 50
rect 1334 16 1360 50
rect 1360 16 1368 50
rect 1406 16 1428 50
rect 1428 16 1440 50
rect 1478 16 1496 50
rect 1496 16 1512 50
rect 1550 16 1564 50
rect 1564 16 1584 50
rect 1622 16 1632 50
rect 1632 16 1656 50
rect 1694 16 1700 50
rect 1700 16 1728 50
rect 1766 16 1768 50
rect 1768 16 1800 50
rect 1838 16 1870 50
rect 1870 16 1872 50
rect 1910 16 1938 50
rect 1938 16 1944 50
rect 1982 16 2006 50
rect 2006 16 2016 50
rect 2054 16 2074 50
rect 2074 16 2088 50
rect 2126 16 2142 50
rect 2142 16 2160 50
rect 2198 16 2210 50
rect 2210 16 2232 50
rect 2270 16 2278 50
rect 2278 16 2304 50
rect 2342 16 2346 50
rect 2346 16 2376 50
rect 2414 16 2448 50
rect 2486 16 2516 50
rect 2516 16 2520 50
rect 2558 16 2584 50
rect 2584 16 2592 50
rect 2630 16 2652 50
rect 2652 16 2664 50
rect 2702 16 2720 50
rect 2720 16 2736 50
rect 2774 16 2788 50
rect 2788 16 2808 50
rect 2846 16 2856 50
rect 2856 16 2880 50
rect 2918 16 2924 50
rect 2924 16 2952 50
rect 2990 16 2992 50
rect 2992 16 3024 50
rect 3062 16 3094 50
rect 3094 16 3096 50
rect 3134 16 3162 50
rect 3162 16 3168 50
rect 3206 16 3230 50
rect 3230 16 3240 50
rect 3278 16 3298 50
rect 3298 16 3312 50
rect 3350 16 3366 50
rect 3366 16 3384 50
rect 3422 16 3434 50
rect 3434 16 3456 50
rect 3494 16 3502 50
rect 3502 16 3528 50
rect 3566 16 3570 50
rect 3570 16 3600 50
rect 3638 16 3672 50
rect 3710 16 3740 50
rect 3740 16 3744 50
rect 3782 16 3808 50
rect 3808 16 3816 50
rect 3854 16 3876 50
rect 3876 16 3888 50
rect 3926 16 3944 50
rect 3944 16 3960 50
rect 3998 16 4012 50
rect 4012 16 4032 50
rect 4070 16 4080 50
rect 4080 16 4104 50
rect 4142 16 4148 50
rect 4148 16 4176 50
rect 4214 16 4216 50
rect 4216 16 4248 50
rect 4286 16 4318 50
rect 4318 16 4320 50
rect 4358 16 4386 50
rect 4386 16 4392 50
<< metal1 >>
rect 0 2331 4498 2338
rect 0 2322 68 2331
rect 120 2322 132 2331
rect 184 2322 292 2331
rect 344 2322 356 2331
rect 408 2322 516 2331
rect 568 2322 580 2331
rect 632 2322 740 2331
rect 0 2288 38 2322
rect 216 2288 254 2322
rect 288 2288 292 2322
rect 432 2288 470 2322
rect 504 2288 516 2322
rect 576 2288 580 2322
rect 648 2288 686 2322
rect 720 2288 740 2322
rect 0 2279 68 2288
rect 120 2279 132 2288
rect 184 2279 292 2288
rect 344 2279 356 2288
rect 408 2279 516 2288
rect 568 2279 580 2288
rect 632 2279 740 2288
rect 792 2279 804 2331
rect 856 2322 964 2331
rect 864 2288 902 2322
rect 936 2288 964 2322
rect 856 2279 964 2288
rect 1016 2279 1028 2331
rect 1080 2322 1188 2331
rect 1080 2288 1118 2322
rect 1152 2288 1188 2322
rect 1080 2279 1188 2288
rect 1240 2279 1252 2331
rect 1304 2322 1412 2331
rect 1304 2288 1334 2322
rect 1368 2288 1406 2322
rect 1304 2279 1412 2288
rect 1464 2279 1476 2331
rect 1528 2322 1636 2331
rect 1688 2322 1700 2331
rect 1752 2322 1860 2331
rect 1912 2322 1924 2331
rect 1976 2322 2084 2331
rect 2136 2322 2148 2331
rect 2200 2322 2308 2331
rect 2360 2322 2372 2331
rect 2424 2322 2532 2331
rect 2584 2322 2596 2331
rect 2648 2322 2756 2331
rect 1528 2288 1550 2322
rect 1584 2288 1622 2322
rect 1688 2288 1694 2322
rect 1752 2288 1766 2322
rect 1800 2288 1838 2322
rect 1976 2288 1982 2322
rect 2016 2288 2054 2322
rect 2232 2288 2270 2322
rect 2304 2288 2308 2322
rect 2448 2288 2486 2322
rect 2520 2288 2532 2322
rect 2592 2288 2596 2322
rect 2664 2288 2702 2322
rect 2736 2288 2756 2322
rect 1528 2279 1636 2288
rect 1688 2279 1700 2288
rect 1752 2279 1860 2288
rect 1912 2279 1924 2288
rect 1976 2279 2084 2288
rect 2136 2279 2148 2288
rect 2200 2279 2308 2288
rect 2360 2279 2372 2288
rect 2424 2279 2532 2288
rect 2584 2279 2596 2288
rect 2648 2279 2756 2288
rect 2808 2279 2820 2331
rect 2872 2322 2980 2331
rect 2880 2288 2918 2322
rect 2952 2288 2980 2322
rect 2872 2279 2980 2288
rect 3032 2279 3044 2331
rect 3096 2322 3204 2331
rect 3096 2288 3134 2322
rect 3168 2288 3204 2322
rect 3096 2279 3204 2288
rect 3256 2279 3268 2331
rect 3320 2322 3428 2331
rect 3320 2288 3350 2322
rect 3384 2288 3422 2322
rect 3320 2279 3428 2288
rect 3480 2279 3492 2331
rect 3544 2322 3652 2331
rect 3704 2322 3716 2331
rect 3768 2322 3876 2331
rect 3928 2322 3940 2331
rect 3992 2322 4100 2331
rect 4152 2322 4164 2331
rect 4216 2322 4324 2331
rect 4376 2322 4388 2331
rect 3544 2288 3566 2322
rect 3600 2288 3638 2322
rect 3704 2288 3710 2322
rect 3768 2288 3782 2322
rect 3816 2288 3854 2322
rect 3992 2288 3998 2322
rect 4032 2288 4070 2322
rect 4248 2288 4286 2322
rect 4320 2288 4324 2322
rect 3544 2279 3652 2288
rect 3704 2279 3716 2288
rect 3768 2279 3876 2288
rect 3928 2279 3940 2288
rect 3992 2279 4100 2288
rect 4152 2279 4164 2288
rect 4216 2279 4324 2288
rect 4376 2279 4388 2288
rect 4440 2279 4498 2331
rect 0 2272 4498 2279
rect 0 94 28 2272
rect 56 66 84 2244
rect 112 94 140 2272
rect 168 66 196 2244
rect 224 94 252 2272
rect 280 66 308 2244
rect 336 94 364 2272
rect 392 66 420 2244
rect 448 94 476 2272
rect 504 66 532 2244
rect 560 94 588 2272
rect 616 66 644 2244
rect 672 94 700 2272
rect 728 66 756 2244
rect 784 94 812 2272
rect 840 66 868 2244
rect 896 94 924 2272
rect 952 66 980 2244
rect 1008 94 1036 2272
rect 1064 66 1092 2244
rect 1120 94 1148 2272
rect 1176 66 1204 2244
rect 1232 94 1260 2272
rect 1288 66 1316 2244
rect 1344 94 1372 2272
rect 1400 66 1428 2244
rect 1456 94 1484 2272
rect 1512 66 1540 2244
rect 1568 94 1596 2272
rect 1624 66 1652 2244
rect 1680 94 1708 2272
rect 1736 66 1764 2244
rect 1792 94 1820 2272
rect 1848 66 1876 2244
rect 1904 94 1932 2272
rect 1960 66 1988 2244
rect 2016 94 2044 2272
rect 2072 66 2100 2244
rect 2128 94 2156 2272
rect 2184 66 2212 2244
rect 2240 94 2268 2272
rect 2296 66 2324 2244
rect 2352 94 2380 2272
rect 2408 66 2436 2244
rect 2464 94 2492 2272
rect 2520 66 2548 2244
rect 2576 94 2604 2272
rect 2632 66 2660 2244
rect 2688 94 2716 2272
rect 2744 66 2772 2244
rect 2800 94 2828 2272
rect 2856 66 2884 2244
rect 2912 94 2940 2272
rect 2968 66 2996 2244
rect 3024 94 3052 2272
rect 3080 66 3108 2244
rect 3136 94 3164 2272
rect 3192 66 3220 2244
rect 3248 94 3276 2272
rect 3304 66 3332 2244
rect 3360 94 3388 2272
rect 3416 66 3444 2244
rect 3472 94 3500 2272
rect 3528 66 3556 2244
rect 3584 94 3612 2272
rect 3640 66 3668 2244
rect 3696 94 3724 2272
rect 3752 66 3780 2244
rect 3808 94 3836 2272
rect 3864 66 3892 2244
rect 3920 94 3948 2272
rect 3976 66 4004 2244
rect 4032 94 4060 2272
rect 4088 66 4116 2244
rect 4144 94 4172 2272
rect 4200 66 4228 2244
rect 4256 94 4284 2272
rect 4312 66 4340 2244
rect 4368 94 4396 2272
rect 4424 66 4498 2244
rect 0 59 4498 66
rect 0 7 24 59
rect 76 7 88 59
rect 140 50 236 59
rect 144 16 182 50
rect 216 16 236 50
rect 140 7 236 16
rect 288 7 300 59
rect 352 50 460 59
rect 360 16 398 50
rect 432 16 460 50
rect 352 7 460 16
rect 512 7 524 59
rect 576 50 684 59
rect 576 16 614 50
rect 648 16 684 50
rect 576 7 684 16
rect 736 7 748 59
rect 800 50 908 59
rect 800 16 830 50
rect 864 16 902 50
rect 800 7 908 16
rect 960 7 972 59
rect 1024 50 1132 59
rect 1184 50 1196 59
rect 1248 50 1356 59
rect 1408 50 1420 59
rect 1472 50 1580 59
rect 1632 50 1644 59
rect 1696 50 1804 59
rect 1856 50 1868 59
rect 1920 50 2028 59
rect 2080 50 2092 59
rect 2144 50 2252 59
rect 1024 16 1046 50
rect 1080 16 1118 50
rect 1184 16 1190 50
rect 1248 16 1262 50
rect 1296 16 1334 50
rect 1472 16 1478 50
rect 1512 16 1550 50
rect 1728 16 1766 50
rect 1800 16 1804 50
rect 1944 16 1982 50
rect 2016 16 2028 50
rect 2088 16 2092 50
rect 2160 16 2198 50
rect 2232 16 2252 50
rect 1024 7 1132 16
rect 1184 7 1196 16
rect 1248 7 1356 16
rect 1408 7 1420 16
rect 1472 7 1580 16
rect 1632 7 1644 16
rect 1696 7 1804 16
rect 1856 7 1868 16
rect 1920 7 2028 16
rect 2080 7 2092 16
rect 2144 7 2252 16
rect 2304 7 2316 59
rect 2368 50 2476 59
rect 2376 16 2414 50
rect 2448 16 2476 50
rect 2368 7 2476 16
rect 2528 7 2540 59
rect 2592 50 2700 59
rect 2592 16 2630 50
rect 2664 16 2700 50
rect 2592 7 2700 16
rect 2752 7 2764 59
rect 2816 50 2924 59
rect 2816 16 2846 50
rect 2880 16 2918 50
rect 2816 7 2924 16
rect 2976 7 2988 59
rect 3040 50 3148 59
rect 3200 50 3212 59
rect 3264 50 3372 59
rect 3424 50 3436 59
rect 3488 50 3596 59
rect 3648 50 3660 59
rect 3712 50 3820 59
rect 3872 50 3884 59
rect 3936 50 4044 59
rect 4096 50 4108 59
rect 4160 50 4268 59
rect 3040 16 3062 50
rect 3096 16 3134 50
rect 3200 16 3206 50
rect 3264 16 3278 50
rect 3312 16 3350 50
rect 3488 16 3494 50
rect 3528 16 3566 50
rect 3744 16 3782 50
rect 3816 16 3820 50
rect 3960 16 3998 50
rect 4032 16 4044 50
rect 4104 16 4108 50
rect 4176 16 4214 50
rect 4248 16 4268 50
rect 3040 7 3148 16
rect 3200 7 3212 16
rect 3264 7 3372 16
rect 3424 7 3436 16
rect 3488 7 3596 16
rect 3648 7 3660 16
rect 3712 7 3820 16
rect 3872 7 3884 16
rect 3936 7 4044 16
rect 4096 7 4108 16
rect 4160 7 4268 16
rect 4320 7 4332 59
rect 4384 50 4498 59
rect 4392 16 4498 50
rect 4384 7 4498 16
rect 0 0 4498 7
<< via1 >>
rect 68 2322 120 2331
rect 132 2322 184 2331
rect 292 2322 344 2331
rect 356 2322 408 2331
rect 516 2322 568 2331
rect 580 2322 632 2331
rect 740 2322 792 2331
rect 68 2288 72 2322
rect 72 2288 110 2322
rect 110 2288 120 2322
rect 132 2288 144 2322
rect 144 2288 182 2322
rect 182 2288 184 2322
rect 292 2288 326 2322
rect 326 2288 344 2322
rect 356 2288 360 2322
rect 360 2288 398 2322
rect 398 2288 408 2322
rect 516 2288 542 2322
rect 542 2288 568 2322
rect 580 2288 614 2322
rect 614 2288 632 2322
rect 740 2288 758 2322
rect 758 2288 792 2322
rect 68 2279 120 2288
rect 132 2279 184 2288
rect 292 2279 344 2288
rect 356 2279 408 2288
rect 516 2279 568 2288
rect 580 2279 632 2288
rect 740 2279 792 2288
rect 804 2322 856 2331
rect 964 2322 1016 2331
rect 804 2288 830 2322
rect 830 2288 856 2322
rect 964 2288 974 2322
rect 974 2288 1008 2322
rect 1008 2288 1016 2322
rect 804 2279 856 2288
rect 964 2279 1016 2288
rect 1028 2322 1080 2331
rect 1188 2322 1240 2331
rect 1028 2288 1046 2322
rect 1046 2288 1080 2322
rect 1188 2288 1190 2322
rect 1190 2288 1224 2322
rect 1224 2288 1240 2322
rect 1028 2279 1080 2288
rect 1188 2279 1240 2288
rect 1252 2322 1304 2331
rect 1412 2322 1464 2331
rect 1252 2288 1262 2322
rect 1262 2288 1296 2322
rect 1296 2288 1304 2322
rect 1412 2288 1440 2322
rect 1440 2288 1464 2322
rect 1252 2279 1304 2288
rect 1412 2279 1464 2288
rect 1476 2322 1528 2331
rect 1636 2322 1688 2331
rect 1700 2322 1752 2331
rect 1860 2322 1912 2331
rect 1924 2322 1976 2331
rect 2084 2322 2136 2331
rect 2148 2322 2200 2331
rect 2308 2322 2360 2331
rect 2372 2322 2424 2331
rect 2532 2322 2584 2331
rect 2596 2322 2648 2331
rect 2756 2322 2808 2331
rect 1476 2288 1478 2322
rect 1478 2288 1512 2322
rect 1512 2288 1528 2322
rect 1636 2288 1656 2322
rect 1656 2288 1688 2322
rect 1700 2288 1728 2322
rect 1728 2288 1752 2322
rect 1860 2288 1872 2322
rect 1872 2288 1910 2322
rect 1910 2288 1912 2322
rect 1924 2288 1944 2322
rect 1944 2288 1976 2322
rect 2084 2288 2088 2322
rect 2088 2288 2126 2322
rect 2126 2288 2136 2322
rect 2148 2288 2160 2322
rect 2160 2288 2198 2322
rect 2198 2288 2200 2322
rect 2308 2288 2342 2322
rect 2342 2288 2360 2322
rect 2372 2288 2376 2322
rect 2376 2288 2414 2322
rect 2414 2288 2424 2322
rect 2532 2288 2558 2322
rect 2558 2288 2584 2322
rect 2596 2288 2630 2322
rect 2630 2288 2648 2322
rect 2756 2288 2774 2322
rect 2774 2288 2808 2322
rect 1476 2279 1528 2288
rect 1636 2279 1688 2288
rect 1700 2279 1752 2288
rect 1860 2279 1912 2288
rect 1924 2279 1976 2288
rect 2084 2279 2136 2288
rect 2148 2279 2200 2288
rect 2308 2279 2360 2288
rect 2372 2279 2424 2288
rect 2532 2279 2584 2288
rect 2596 2279 2648 2288
rect 2756 2279 2808 2288
rect 2820 2322 2872 2331
rect 2980 2322 3032 2331
rect 2820 2288 2846 2322
rect 2846 2288 2872 2322
rect 2980 2288 2990 2322
rect 2990 2288 3024 2322
rect 3024 2288 3032 2322
rect 2820 2279 2872 2288
rect 2980 2279 3032 2288
rect 3044 2322 3096 2331
rect 3204 2322 3256 2331
rect 3044 2288 3062 2322
rect 3062 2288 3096 2322
rect 3204 2288 3206 2322
rect 3206 2288 3240 2322
rect 3240 2288 3256 2322
rect 3044 2279 3096 2288
rect 3204 2279 3256 2288
rect 3268 2322 3320 2331
rect 3428 2322 3480 2331
rect 3268 2288 3278 2322
rect 3278 2288 3312 2322
rect 3312 2288 3320 2322
rect 3428 2288 3456 2322
rect 3456 2288 3480 2322
rect 3268 2279 3320 2288
rect 3428 2279 3480 2288
rect 3492 2322 3544 2331
rect 3652 2322 3704 2331
rect 3716 2322 3768 2331
rect 3876 2322 3928 2331
rect 3940 2322 3992 2331
rect 4100 2322 4152 2331
rect 4164 2322 4216 2331
rect 4324 2322 4376 2331
rect 4388 2322 4440 2331
rect 3492 2288 3494 2322
rect 3494 2288 3528 2322
rect 3528 2288 3544 2322
rect 3652 2288 3672 2322
rect 3672 2288 3704 2322
rect 3716 2288 3744 2322
rect 3744 2288 3768 2322
rect 3876 2288 3888 2322
rect 3888 2288 3926 2322
rect 3926 2288 3928 2322
rect 3940 2288 3960 2322
rect 3960 2288 3992 2322
rect 4100 2288 4104 2322
rect 4104 2288 4142 2322
rect 4142 2288 4152 2322
rect 4164 2288 4176 2322
rect 4176 2288 4214 2322
rect 4214 2288 4216 2322
rect 4324 2288 4358 2322
rect 4358 2288 4376 2322
rect 4388 2288 4392 2322
rect 4392 2288 4440 2322
rect 3492 2279 3544 2288
rect 3652 2279 3704 2288
rect 3716 2279 3768 2288
rect 3876 2279 3928 2288
rect 3940 2279 3992 2288
rect 4100 2279 4152 2288
rect 4164 2279 4216 2288
rect 4324 2279 4376 2288
rect 4388 2279 4440 2288
rect 24 50 76 59
rect 24 16 38 50
rect 38 16 72 50
rect 72 16 76 50
rect 24 7 76 16
rect 88 50 140 59
rect 236 50 288 59
rect 88 16 110 50
rect 110 16 140 50
rect 236 16 254 50
rect 254 16 288 50
rect 88 7 140 16
rect 236 7 288 16
rect 300 50 352 59
rect 460 50 512 59
rect 300 16 326 50
rect 326 16 352 50
rect 460 16 470 50
rect 470 16 504 50
rect 504 16 512 50
rect 300 7 352 16
rect 460 7 512 16
rect 524 50 576 59
rect 684 50 736 59
rect 524 16 542 50
rect 542 16 576 50
rect 684 16 686 50
rect 686 16 720 50
rect 720 16 736 50
rect 524 7 576 16
rect 684 7 736 16
rect 748 50 800 59
rect 908 50 960 59
rect 748 16 758 50
rect 758 16 792 50
rect 792 16 800 50
rect 908 16 936 50
rect 936 16 960 50
rect 748 7 800 16
rect 908 7 960 16
rect 972 50 1024 59
rect 1132 50 1184 59
rect 1196 50 1248 59
rect 1356 50 1408 59
rect 1420 50 1472 59
rect 1580 50 1632 59
rect 1644 50 1696 59
rect 1804 50 1856 59
rect 1868 50 1920 59
rect 2028 50 2080 59
rect 2092 50 2144 59
rect 2252 50 2304 59
rect 972 16 974 50
rect 974 16 1008 50
rect 1008 16 1024 50
rect 1132 16 1152 50
rect 1152 16 1184 50
rect 1196 16 1224 50
rect 1224 16 1248 50
rect 1356 16 1368 50
rect 1368 16 1406 50
rect 1406 16 1408 50
rect 1420 16 1440 50
rect 1440 16 1472 50
rect 1580 16 1584 50
rect 1584 16 1622 50
rect 1622 16 1632 50
rect 1644 16 1656 50
rect 1656 16 1694 50
rect 1694 16 1696 50
rect 1804 16 1838 50
rect 1838 16 1856 50
rect 1868 16 1872 50
rect 1872 16 1910 50
rect 1910 16 1920 50
rect 2028 16 2054 50
rect 2054 16 2080 50
rect 2092 16 2126 50
rect 2126 16 2144 50
rect 2252 16 2270 50
rect 2270 16 2304 50
rect 972 7 1024 16
rect 1132 7 1184 16
rect 1196 7 1248 16
rect 1356 7 1408 16
rect 1420 7 1472 16
rect 1580 7 1632 16
rect 1644 7 1696 16
rect 1804 7 1856 16
rect 1868 7 1920 16
rect 2028 7 2080 16
rect 2092 7 2144 16
rect 2252 7 2304 16
rect 2316 50 2368 59
rect 2476 50 2528 59
rect 2316 16 2342 50
rect 2342 16 2368 50
rect 2476 16 2486 50
rect 2486 16 2520 50
rect 2520 16 2528 50
rect 2316 7 2368 16
rect 2476 7 2528 16
rect 2540 50 2592 59
rect 2700 50 2752 59
rect 2540 16 2558 50
rect 2558 16 2592 50
rect 2700 16 2702 50
rect 2702 16 2736 50
rect 2736 16 2752 50
rect 2540 7 2592 16
rect 2700 7 2752 16
rect 2764 50 2816 59
rect 2924 50 2976 59
rect 2764 16 2774 50
rect 2774 16 2808 50
rect 2808 16 2816 50
rect 2924 16 2952 50
rect 2952 16 2976 50
rect 2764 7 2816 16
rect 2924 7 2976 16
rect 2988 50 3040 59
rect 3148 50 3200 59
rect 3212 50 3264 59
rect 3372 50 3424 59
rect 3436 50 3488 59
rect 3596 50 3648 59
rect 3660 50 3712 59
rect 3820 50 3872 59
rect 3884 50 3936 59
rect 4044 50 4096 59
rect 4108 50 4160 59
rect 4268 50 4320 59
rect 2988 16 2990 50
rect 2990 16 3024 50
rect 3024 16 3040 50
rect 3148 16 3168 50
rect 3168 16 3200 50
rect 3212 16 3240 50
rect 3240 16 3264 50
rect 3372 16 3384 50
rect 3384 16 3422 50
rect 3422 16 3424 50
rect 3436 16 3456 50
rect 3456 16 3488 50
rect 3596 16 3600 50
rect 3600 16 3638 50
rect 3638 16 3648 50
rect 3660 16 3672 50
rect 3672 16 3710 50
rect 3710 16 3712 50
rect 3820 16 3854 50
rect 3854 16 3872 50
rect 3884 16 3888 50
rect 3888 16 3926 50
rect 3926 16 3936 50
rect 4044 16 4070 50
rect 4070 16 4096 50
rect 4108 16 4142 50
rect 4142 16 4160 50
rect 4268 16 4286 50
rect 4286 16 4320 50
rect 2988 7 3040 16
rect 3148 7 3200 16
rect 3212 7 3264 16
rect 3372 7 3424 16
rect 3436 7 3488 16
rect 3596 7 3648 16
rect 3660 7 3712 16
rect 3820 7 3872 16
rect 3884 7 3936 16
rect 4044 7 4096 16
rect 4108 7 4160 16
rect 4268 7 4320 16
rect 4332 50 4384 59
rect 4332 16 4358 50
rect 4358 16 4384 50
rect 4332 7 4384 16
<< metal2 >>
rect 0 66 28 2338
rect 56 2333 196 2338
rect 56 2331 98 2333
rect 154 2331 196 2333
rect 56 2279 68 2331
rect 184 2279 196 2331
rect 56 2277 98 2279
rect 154 2277 196 2279
rect 56 2272 196 2277
rect 56 94 84 2272
rect 112 66 140 2244
rect 0 61 140 66
rect 0 59 42 61
rect 98 59 140 61
rect 0 7 24 59
rect 0 5 42 7
rect 98 5 140 7
rect 0 0 140 5
rect 168 0 196 2272
rect 224 66 252 2338
rect 280 2333 420 2338
rect 280 2331 322 2333
rect 378 2331 420 2333
rect 280 2279 292 2331
rect 408 2279 420 2331
rect 280 2277 322 2279
rect 378 2277 420 2279
rect 280 2272 420 2277
rect 280 94 308 2272
rect 336 66 364 2244
rect 224 61 364 66
rect 224 59 266 61
rect 322 59 364 61
rect 224 7 236 59
rect 352 7 364 59
rect 224 5 266 7
rect 322 5 364 7
rect 224 0 364 5
rect 392 0 420 2272
rect 448 66 476 2338
rect 504 2333 644 2338
rect 504 2331 546 2333
rect 602 2331 644 2333
rect 504 2279 516 2331
rect 632 2279 644 2331
rect 504 2277 546 2279
rect 602 2277 644 2279
rect 504 2272 644 2277
rect 504 94 532 2272
rect 560 66 588 2244
rect 448 61 588 66
rect 448 59 490 61
rect 546 59 588 61
rect 448 7 460 59
rect 576 7 588 59
rect 448 5 490 7
rect 546 5 588 7
rect 448 0 588 5
rect 616 0 644 2272
rect 672 66 700 2338
rect 728 2333 868 2338
rect 728 2331 770 2333
rect 826 2331 868 2333
rect 728 2279 740 2331
rect 856 2279 868 2331
rect 728 2277 770 2279
rect 826 2277 868 2279
rect 728 2272 868 2277
rect 728 94 756 2272
rect 784 66 812 2244
rect 672 61 812 66
rect 672 59 714 61
rect 770 59 812 61
rect 672 7 684 59
rect 800 7 812 59
rect 672 5 714 7
rect 770 5 812 7
rect 672 0 812 5
rect 840 0 868 2272
rect 896 66 924 2338
rect 952 2333 1092 2338
rect 952 2331 994 2333
rect 1050 2331 1092 2333
rect 952 2279 964 2331
rect 1080 2279 1092 2331
rect 952 2277 994 2279
rect 1050 2277 1092 2279
rect 952 2272 1092 2277
rect 952 94 980 2272
rect 1008 66 1036 2244
rect 896 61 1036 66
rect 896 59 938 61
rect 994 59 1036 61
rect 896 7 908 59
rect 1024 7 1036 59
rect 896 5 938 7
rect 994 5 1036 7
rect 896 0 1036 5
rect 1064 0 1092 2272
rect 1120 66 1148 2338
rect 1176 2333 1316 2338
rect 1176 2331 1218 2333
rect 1274 2331 1316 2333
rect 1176 2279 1188 2331
rect 1304 2279 1316 2331
rect 1176 2277 1218 2279
rect 1274 2277 1316 2279
rect 1176 2272 1316 2277
rect 1176 94 1204 2272
rect 1232 66 1260 2244
rect 1120 61 1260 66
rect 1120 59 1162 61
rect 1218 59 1260 61
rect 1120 7 1132 59
rect 1248 7 1260 59
rect 1120 5 1162 7
rect 1218 5 1260 7
rect 1120 0 1260 5
rect 1288 0 1316 2272
rect 1344 66 1372 2338
rect 1400 2333 1540 2338
rect 1400 2331 1442 2333
rect 1498 2331 1540 2333
rect 1400 2279 1412 2331
rect 1528 2279 1540 2331
rect 1400 2277 1442 2279
rect 1498 2277 1540 2279
rect 1400 2272 1540 2277
rect 1400 94 1428 2272
rect 1456 66 1484 2244
rect 1344 61 1484 66
rect 1344 59 1386 61
rect 1442 59 1484 61
rect 1344 7 1356 59
rect 1472 7 1484 59
rect 1344 5 1386 7
rect 1442 5 1484 7
rect 1344 0 1484 5
rect 1512 0 1540 2272
rect 1568 66 1596 2338
rect 1624 2333 1764 2338
rect 1624 2331 1666 2333
rect 1722 2331 1764 2333
rect 1624 2279 1636 2331
rect 1752 2279 1764 2331
rect 1624 2277 1666 2279
rect 1722 2277 1764 2279
rect 1624 2272 1764 2277
rect 1624 94 1652 2272
rect 1680 66 1708 2244
rect 1568 61 1708 66
rect 1568 59 1610 61
rect 1666 59 1708 61
rect 1568 7 1580 59
rect 1696 7 1708 59
rect 1568 5 1610 7
rect 1666 5 1708 7
rect 1568 0 1708 5
rect 1736 0 1764 2272
rect 1792 66 1820 2338
rect 1848 2333 1988 2338
rect 1848 2331 1890 2333
rect 1946 2331 1988 2333
rect 1848 2279 1860 2331
rect 1976 2279 1988 2331
rect 1848 2277 1890 2279
rect 1946 2277 1988 2279
rect 1848 2272 1988 2277
rect 1848 94 1876 2272
rect 1904 66 1932 2244
rect 1792 61 1932 66
rect 1792 59 1834 61
rect 1890 59 1932 61
rect 1792 7 1804 59
rect 1920 7 1932 59
rect 1792 5 1834 7
rect 1890 5 1932 7
rect 1792 0 1932 5
rect 1960 0 1988 2272
rect 2016 66 2044 2338
rect 2072 2333 2212 2338
rect 2072 2331 2114 2333
rect 2170 2331 2212 2333
rect 2072 2279 2084 2331
rect 2200 2279 2212 2331
rect 2072 2277 2114 2279
rect 2170 2277 2212 2279
rect 2072 2272 2212 2277
rect 2072 94 2100 2272
rect 2128 66 2156 2244
rect 2016 61 2156 66
rect 2016 59 2058 61
rect 2114 59 2156 61
rect 2016 7 2028 59
rect 2144 7 2156 59
rect 2016 5 2058 7
rect 2114 5 2156 7
rect 2016 0 2156 5
rect 2184 0 2212 2272
rect 2240 66 2268 2338
rect 2296 2333 2436 2338
rect 2296 2331 2338 2333
rect 2394 2331 2436 2333
rect 2296 2279 2308 2331
rect 2424 2279 2436 2331
rect 2296 2277 2338 2279
rect 2394 2277 2436 2279
rect 2296 2272 2436 2277
rect 2296 94 2324 2272
rect 2352 66 2380 2244
rect 2240 61 2380 66
rect 2240 59 2282 61
rect 2338 59 2380 61
rect 2240 7 2252 59
rect 2368 7 2380 59
rect 2240 5 2282 7
rect 2338 5 2380 7
rect 2240 0 2380 5
rect 2408 0 2436 2272
rect 2464 66 2492 2338
rect 2520 2333 2660 2338
rect 2520 2331 2562 2333
rect 2618 2331 2660 2333
rect 2520 2279 2532 2331
rect 2648 2279 2660 2331
rect 2520 2277 2562 2279
rect 2618 2277 2660 2279
rect 2520 2272 2660 2277
rect 2520 94 2548 2272
rect 2576 66 2604 2244
rect 2464 61 2604 66
rect 2464 59 2506 61
rect 2562 59 2604 61
rect 2464 7 2476 59
rect 2592 7 2604 59
rect 2464 5 2506 7
rect 2562 5 2604 7
rect 2464 0 2604 5
rect 2632 0 2660 2272
rect 2688 66 2716 2338
rect 2744 2333 2884 2338
rect 2744 2331 2786 2333
rect 2842 2331 2884 2333
rect 2744 2279 2756 2331
rect 2872 2279 2884 2331
rect 2744 2277 2786 2279
rect 2842 2277 2884 2279
rect 2744 2272 2884 2277
rect 2744 94 2772 2272
rect 2800 66 2828 2244
rect 2688 61 2828 66
rect 2688 59 2730 61
rect 2786 59 2828 61
rect 2688 7 2700 59
rect 2816 7 2828 59
rect 2688 5 2730 7
rect 2786 5 2828 7
rect 2688 0 2828 5
rect 2856 0 2884 2272
rect 2912 66 2940 2338
rect 2968 2333 3108 2338
rect 2968 2331 3010 2333
rect 3066 2331 3108 2333
rect 2968 2279 2980 2331
rect 3096 2279 3108 2331
rect 2968 2277 3010 2279
rect 3066 2277 3108 2279
rect 2968 2272 3108 2277
rect 2968 94 2996 2272
rect 3024 66 3052 2244
rect 2912 61 3052 66
rect 2912 59 2954 61
rect 3010 59 3052 61
rect 2912 7 2924 59
rect 3040 7 3052 59
rect 2912 5 2954 7
rect 3010 5 3052 7
rect 2912 0 3052 5
rect 3080 0 3108 2272
rect 3136 66 3164 2338
rect 3192 2333 3332 2338
rect 3192 2331 3234 2333
rect 3290 2331 3332 2333
rect 3192 2279 3204 2331
rect 3320 2279 3332 2331
rect 3192 2277 3234 2279
rect 3290 2277 3332 2279
rect 3192 2272 3332 2277
rect 3192 94 3220 2272
rect 3248 66 3276 2244
rect 3136 61 3276 66
rect 3136 59 3178 61
rect 3234 59 3276 61
rect 3136 7 3148 59
rect 3264 7 3276 59
rect 3136 5 3178 7
rect 3234 5 3276 7
rect 3136 0 3276 5
rect 3304 0 3332 2272
rect 3360 66 3388 2338
rect 3416 2333 3556 2338
rect 3416 2331 3458 2333
rect 3514 2331 3556 2333
rect 3416 2279 3428 2331
rect 3544 2279 3556 2331
rect 3416 2277 3458 2279
rect 3514 2277 3556 2279
rect 3416 2272 3556 2277
rect 3416 94 3444 2272
rect 3472 66 3500 2244
rect 3360 61 3500 66
rect 3360 59 3402 61
rect 3458 59 3500 61
rect 3360 7 3372 59
rect 3488 7 3500 59
rect 3360 5 3402 7
rect 3458 5 3500 7
rect 3360 0 3500 5
rect 3528 0 3556 2272
rect 3584 66 3612 2338
rect 3640 2333 3780 2338
rect 3640 2331 3682 2333
rect 3738 2331 3780 2333
rect 3640 2279 3652 2331
rect 3768 2279 3780 2331
rect 3640 2277 3682 2279
rect 3738 2277 3780 2279
rect 3640 2272 3780 2277
rect 3640 94 3668 2272
rect 3696 66 3724 2244
rect 3584 61 3724 66
rect 3584 59 3626 61
rect 3682 59 3724 61
rect 3584 7 3596 59
rect 3712 7 3724 59
rect 3584 5 3626 7
rect 3682 5 3724 7
rect 3584 0 3724 5
rect 3752 0 3780 2272
rect 3808 66 3836 2338
rect 3864 2333 4004 2338
rect 3864 2331 3906 2333
rect 3962 2331 4004 2333
rect 3864 2279 3876 2331
rect 3992 2279 4004 2331
rect 3864 2277 3906 2279
rect 3962 2277 4004 2279
rect 3864 2272 4004 2277
rect 3864 94 3892 2272
rect 3920 66 3948 2244
rect 3808 61 3948 66
rect 3808 59 3850 61
rect 3906 59 3948 61
rect 3808 7 3820 59
rect 3936 7 3948 59
rect 3808 5 3850 7
rect 3906 5 3948 7
rect 3808 0 3948 5
rect 3976 0 4004 2272
rect 4032 66 4060 2338
rect 4088 2333 4498 2338
rect 4088 2331 4130 2333
rect 4186 2331 4498 2333
rect 4088 2279 4100 2331
rect 4216 2279 4324 2331
rect 4376 2279 4388 2331
rect 4440 2279 4498 2331
rect 4088 2277 4130 2279
rect 4186 2277 4498 2279
rect 4088 2272 4498 2277
rect 4088 94 4116 2272
rect 4144 66 4172 2244
rect 4032 61 4172 66
rect 4032 59 4074 61
rect 4130 59 4172 61
rect 4032 7 4044 59
rect 4160 7 4172 59
rect 4032 5 4074 7
rect 4130 5 4172 7
rect 4032 0 4172 5
rect 4200 0 4228 2272
rect 4256 66 4284 2244
rect 4312 94 4340 2272
rect 4368 66 4396 2244
rect 4424 94 4498 2272
rect 4256 61 4498 66
rect 4256 59 4298 61
rect 4354 59 4498 61
rect 4256 7 4268 59
rect 4384 7 4498 59
rect 4256 5 4298 7
rect 4354 5 4498 7
rect 4256 0 4498 5
<< via2 >>
rect 98 2331 154 2333
rect 98 2279 120 2331
rect 120 2279 132 2331
rect 132 2279 154 2331
rect 98 2277 154 2279
rect 42 59 98 61
rect 42 7 76 59
rect 76 7 88 59
rect 88 7 98 59
rect 42 5 98 7
rect 322 2331 378 2333
rect 322 2279 344 2331
rect 344 2279 356 2331
rect 356 2279 378 2331
rect 322 2277 378 2279
rect 266 59 322 61
rect 266 7 288 59
rect 288 7 300 59
rect 300 7 322 59
rect 266 5 322 7
rect 546 2331 602 2333
rect 546 2279 568 2331
rect 568 2279 580 2331
rect 580 2279 602 2331
rect 546 2277 602 2279
rect 490 59 546 61
rect 490 7 512 59
rect 512 7 524 59
rect 524 7 546 59
rect 490 5 546 7
rect 770 2331 826 2333
rect 770 2279 792 2331
rect 792 2279 804 2331
rect 804 2279 826 2331
rect 770 2277 826 2279
rect 714 59 770 61
rect 714 7 736 59
rect 736 7 748 59
rect 748 7 770 59
rect 714 5 770 7
rect 994 2331 1050 2333
rect 994 2279 1016 2331
rect 1016 2279 1028 2331
rect 1028 2279 1050 2331
rect 994 2277 1050 2279
rect 938 59 994 61
rect 938 7 960 59
rect 960 7 972 59
rect 972 7 994 59
rect 938 5 994 7
rect 1218 2331 1274 2333
rect 1218 2279 1240 2331
rect 1240 2279 1252 2331
rect 1252 2279 1274 2331
rect 1218 2277 1274 2279
rect 1162 59 1218 61
rect 1162 7 1184 59
rect 1184 7 1196 59
rect 1196 7 1218 59
rect 1162 5 1218 7
rect 1442 2331 1498 2333
rect 1442 2279 1464 2331
rect 1464 2279 1476 2331
rect 1476 2279 1498 2331
rect 1442 2277 1498 2279
rect 1386 59 1442 61
rect 1386 7 1408 59
rect 1408 7 1420 59
rect 1420 7 1442 59
rect 1386 5 1442 7
rect 1666 2331 1722 2333
rect 1666 2279 1688 2331
rect 1688 2279 1700 2331
rect 1700 2279 1722 2331
rect 1666 2277 1722 2279
rect 1610 59 1666 61
rect 1610 7 1632 59
rect 1632 7 1644 59
rect 1644 7 1666 59
rect 1610 5 1666 7
rect 1890 2331 1946 2333
rect 1890 2279 1912 2331
rect 1912 2279 1924 2331
rect 1924 2279 1946 2331
rect 1890 2277 1946 2279
rect 1834 59 1890 61
rect 1834 7 1856 59
rect 1856 7 1868 59
rect 1868 7 1890 59
rect 1834 5 1890 7
rect 2114 2331 2170 2333
rect 2114 2279 2136 2331
rect 2136 2279 2148 2331
rect 2148 2279 2170 2331
rect 2114 2277 2170 2279
rect 2058 59 2114 61
rect 2058 7 2080 59
rect 2080 7 2092 59
rect 2092 7 2114 59
rect 2058 5 2114 7
rect 2338 2331 2394 2333
rect 2338 2279 2360 2331
rect 2360 2279 2372 2331
rect 2372 2279 2394 2331
rect 2338 2277 2394 2279
rect 2282 59 2338 61
rect 2282 7 2304 59
rect 2304 7 2316 59
rect 2316 7 2338 59
rect 2282 5 2338 7
rect 2562 2331 2618 2333
rect 2562 2279 2584 2331
rect 2584 2279 2596 2331
rect 2596 2279 2618 2331
rect 2562 2277 2618 2279
rect 2506 59 2562 61
rect 2506 7 2528 59
rect 2528 7 2540 59
rect 2540 7 2562 59
rect 2506 5 2562 7
rect 2786 2331 2842 2333
rect 2786 2279 2808 2331
rect 2808 2279 2820 2331
rect 2820 2279 2842 2331
rect 2786 2277 2842 2279
rect 2730 59 2786 61
rect 2730 7 2752 59
rect 2752 7 2764 59
rect 2764 7 2786 59
rect 2730 5 2786 7
rect 3010 2331 3066 2333
rect 3010 2279 3032 2331
rect 3032 2279 3044 2331
rect 3044 2279 3066 2331
rect 3010 2277 3066 2279
rect 2954 59 3010 61
rect 2954 7 2976 59
rect 2976 7 2988 59
rect 2988 7 3010 59
rect 2954 5 3010 7
rect 3234 2331 3290 2333
rect 3234 2279 3256 2331
rect 3256 2279 3268 2331
rect 3268 2279 3290 2331
rect 3234 2277 3290 2279
rect 3178 59 3234 61
rect 3178 7 3200 59
rect 3200 7 3212 59
rect 3212 7 3234 59
rect 3178 5 3234 7
rect 3458 2331 3514 2333
rect 3458 2279 3480 2331
rect 3480 2279 3492 2331
rect 3492 2279 3514 2331
rect 3458 2277 3514 2279
rect 3402 59 3458 61
rect 3402 7 3424 59
rect 3424 7 3436 59
rect 3436 7 3458 59
rect 3402 5 3458 7
rect 3682 2331 3738 2333
rect 3682 2279 3704 2331
rect 3704 2279 3716 2331
rect 3716 2279 3738 2331
rect 3682 2277 3738 2279
rect 3626 59 3682 61
rect 3626 7 3648 59
rect 3648 7 3660 59
rect 3660 7 3682 59
rect 3626 5 3682 7
rect 3906 2331 3962 2333
rect 3906 2279 3928 2331
rect 3928 2279 3940 2331
rect 3940 2279 3962 2331
rect 3906 2277 3962 2279
rect 3850 59 3906 61
rect 3850 7 3872 59
rect 3872 7 3884 59
rect 3884 7 3906 59
rect 3850 5 3906 7
rect 4130 2331 4186 2333
rect 4130 2279 4152 2331
rect 4152 2279 4164 2331
rect 4164 2279 4186 2331
rect 4130 2277 4186 2279
rect 4074 59 4130 61
rect 4074 7 4096 59
rect 4096 7 4108 59
rect 4108 7 4130 59
rect 4074 5 4130 7
rect 4298 59 4354 61
rect 4298 7 4320 59
rect 4320 7 4332 59
rect 4332 7 4354 59
rect 4298 5 4354 7
<< metal3 >>
rect 0 2337 4498 2338
rect 0 2273 28 2337
rect 92 2333 108 2337
rect 92 2277 98 2333
rect 92 2273 108 2277
rect 172 2273 188 2337
rect 252 2273 268 2337
rect 332 2333 348 2337
rect 332 2273 348 2277
rect 412 2273 428 2337
rect 492 2273 508 2337
rect 572 2333 588 2337
rect 572 2273 588 2277
rect 652 2273 668 2337
rect 732 2273 748 2337
rect 812 2333 828 2337
rect 826 2277 828 2333
rect 812 2273 828 2277
rect 892 2273 908 2337
rect 972 2273 988 2337
rect 1052 2273 1068 2337
rect 1132 2273 1148 2337
rect 1212 2333 1228 2337
rect 1212 2277 1218 2333
rect 1212 2273 1228 2277
rect 1292 2273 1308 2337
rect 1372 2273 1388 2337
rect 1452 2333 1468 2337
rect 1452 2273 1468 2277
rect 1532 2273 1548 2337
rect 1612 2273 1628 2337
rect 1692 2333 1708 2337
rect 1692 2273 1708 2277
rect 1772 2273 1788 2337
rect 1852 2273 1868 2337
rect 1932 2333 1948 2337
rect 1946 2277 1948 2333
rect 1932 2273 1948 2277
rect 2012 2273 2028 2337
rect 2092 2273 2108 2337
rect 2172 2273 2188 2337
rect 2252 2273 2268 2337
rect 2332 2333 2348 2337
rect 2332 2277 2338 2333
rect 2332 2273 2348 2277
rect 2412 2273 2428 2337
rect 2492 2273 2508 2337
rect 2572 2333 2588 2337
rect 2572 2273 2588 2277
rect 2652 2273 2668 2337
rect 2732 2273 2748 2337
rect 2812 2333 2828 2337
rect 2812 2273 2828 2277
rect 2892 2273 2908 2337
rect 2972 2273 2988 2337
rect 3052 2333 3068 2337
rect 3066 2277 3068 2333
rect 3052 2273 3068 2277
rect 3132 2273 3148 2337
rect 3212 2273 3228 2337
rect 3292 2273 3308 2337
rect 3372 2273 3388 2337
rect 3452 2333 3468 2337
rect 3452 2277 3458 2333
rect 3452 2273 3468 2277
rect 3532 2273 3548 2337
rect 3612 2273 3628 2337
rect 3692 2333 3708 2337
rect 3692 2273 3708 2277
rect 3772 2273 3788 2337
rect 3852 2273 3868 2337
rect 3932 2333 3948 2337
rect 3932 2273 3948 2277
rect 4012 2273 4028 2337
rect 4092 2273 4108 2337
rect 4172 2333 4188 2337
rect 4186 2277 4188 2333
rect 4172 2273 4188 2277
rect 4252 2273 4268 2337
rect 4332 2273 4348 2337
rect 4412 2273 4498 2337
rect 0 2272 4498 2273
rect 0 126 60 2272
rect 120 66 180 2212
rect 240 126 300 2272
rect 360 66 420 2212
rect 480 126 540 2272
rect 600 66 660 2212
rect 720 126 780 2272
rect 840 66 900 2212
rect 960 126 1020 2272
rect 1080 66 1140 2212
rect 1200 126 1260 2272
rect 1320 66 1380 2212
rect 1440 126 1500 2272
rect 1560 66 1620 2212
rect 1680 126 1740 2272
rect 1800 66 1860 2212
rect 1920 126 1980 2272
rect 2040 66 2100 2212
rect 2160 126 2220 2272
rect 2280 66 2340 2212
rect 2400 126 2460 2272
rect 2520 66 2580 2212
rect 2640 126 2700 2272
rect 2760 66 2820 2212
rect 2880 126 2940 2272
rect 3000 66 3060 2212
rect 3120 126 3180 2272
rect 3240 66 3300 2212
rect 3360 126 3420 2272
rect 3480 66 3540 2212
rect 3600 126 3660 2272
rect 3720 66 3780 2212
rect 3840 126 3900 2272
rect 3960 66 4020 2212
rect 4080 126 4140 2272
rect 4200 66 4260 2212
rect 4320 126 4498 2272
rect 0 65 4498 66
rect 0 1 28 65
rect 92 61 108 65
rect 98 5 108 61
rect 92 1 108 5
rect 172 1 188 65
rect 252 61 268 65
rect 252 5 266 61
rect 252 1 268 5
rect 332 1 348 65
rect 412 1 428 65
rect 492 61 508 65
rect 492 1 508 5
rect 572 1 588 65
rect 652 1 668 65
rect 732 61 748 65
rect 732 1 748 5
rect 812 1 828 65
rect 892 1 908 65
rect 972 61 988 65
rect 972 1 988 5
rect 1052 1 1068 65
rect 1132 1 1148 65
rect 1212 61 1228 65
rect 1218 5 1228 61
rect 1212 1 1228 5
rect 1292 1 1308 65
rect 1372 61 1388 65
rect 1372 5 1386 61
rect 1372 1 1388 5
rect 1452 1 1468 65
rect 1532 1 1548 65
rect 1612 61 1628 65
rect 1612 1 1628 5
rect 1692 1 1708 65
rect 1772 1 1788 65
rect 1852 61 1868 65
rect 1852 1 1868 5
rect 1932 1 1948 65
rect 2012 1 2028 65
rect 2092 61 2108 65
rect 2092 1 2108 5
rect 2172 1 2188 65
rect 2252 1 2268 65
rect 2332 61 2348 65
rect 2338 5 2348 61
rect 2332 1 2348 5
rect 2412 1 2428 65
rect 2492 61 2508 65
rect 2492 5 2506 61
rect 2492 1 2508 5
rect 2572 1 2588 65
rect 2652 1 2668 65
rect 2732 61 2748 65
rect 2732 1 2748 5
rect 2812 1 2828 65
rect 2892 1 2908 65
rect 2972 61 2988 65
rect 2972 1 2988 5
rect 3052 1 3068 65
rect 3132 1 3148 65
rect 3212 61 3228 65
rect 3212 1 3228 5
rect 3292 1 3308 65
rect 3372 1 3388 65
rect 3452 61 3468 65
rect 3458 5 3468 61
rect 3452 1 3468 5
rect 3532 1 3548 65
rect 3612 61 3628 65
rect 3612 5 3626 61
rect 3612 1 3628 5
rect 3692 1 3708 65
rect 3772 1 3788 65
rect 3852 61 3868 65
rect 3852 1 3868 5
rect 3932 1 3948 65
rect 4012 1 4028 65
rect 4092 61 4108 65
rect 4092 1 4108 5
rect 4172 1 4188 65
rect 4252 1 4268 65
rect 4332 61 4348 65
rect 4332 1 4348 5
rect 4412 1 4498 65
rect 0 0 4498 1
<< via3 >>
rect 28 2273 92 2337
rect 108 2333 172 2337
rect 108 2277 154 2333
rect 154 2277 172 2333
rect 108 2273 172 2277
rect 188 2273 252 2337
rect 268 2333 332 2337
rect 348 2333 412 2337
rect 268 2277 322 2333
rect 322 2277 332 2333
rect 348 2277 378 2333
rect 378 2277 412 2333
rect 268 2273 332 2277
rect 348 2273 412 2277
rect 428 2273 492 2337
rect 508 2333 572 2337
rect 588 2333 652 2337
rect 508 2277 546 2333
rect 546 2277 572 2333
rect 588 2277 602 2333
rect 602 2277 652 2333
rect 508 2273 572 2277
rect 588 2273 652 2277
rect 668 2273 732 2337
rect 748 2333 812 2337
rect 748 2277 770 2333
rect 770 2277 812 2333
rect 748 2273 812 2277
rect 828 2273 892 2337
rect 908 2273 972 2337
rect 988 2333 1052 2337
rect 988 2277 994 2333
rect 994 2277 1050 2333
rect 1050 2277 1052 2333
rect 988 2273 1052 2277
rect 1068 2273 1132 2337
rect 1148 2273 1212 2337
rect 1228 2333 1292 2337
rect 1228 2277 1274 2333
rect 1274 2277 1292 2333
rect 1228 2273 1292 2277
rect 1308 2273 1372 2337
rect 1388 2333 1452 2337
rect 1468 2333 1532 2337
rect 1388 2277 1442 2333
rect 1442 2277 1452 2333
rect 1468 2277 1498 2333
rect 1498 2277 1532 2333
rect 1388 2273 1452 2277
rect 1468 2273 1532 2277
rect 1548 2273 1612 2337
rect 1628 2333 1692 2337
rect 1708 2333 1772 2337
rect 1628 2277 1666 2333
rect 1666 2277 1692 2333
rect 1708 2277 1722 2333
rect 1722 2277 1772 2333
rect 1628 2273 1692 2277
rect 1708 2273 1772 2277
rect 1788 2273 1852 2337
rect 1868 2333 1932 2337
rect 1868 2277 1890 2333
rect 1890 2277 1932 2333
rect 1868 2273 1932 2277
rect 1948 2273 2012 2337
rect 2028 2273 2092 2337
rect 2108 2333 2172 2337
rect 2108 2277 2114 2333
rect 2114 2277 2170 2333
rect 2170 2277 2172 2333
rect 2108 2273 2172 2277
rect 2188 2273 2252 2337
rect 2268 2273 2332 2337
rect 2348 2333 2412 2337
rect 2348 2277 2394 2333
rect 2394 2277 2412 2333
rect 2348 2273 2412 2277
rect 2428 2273 2492 2337
rect 2508 2333 2572 2337
rect 2588 2333 2652 2337
rect 2508 2277 2562 2333
rect 2562 2277 2572 2333
rect 2588 2277 2618 2333
rect 2618 2277 2652 2333
rect 2508 2273 2572 2277
rect 2588 2273 2652 2277
rect 2668 2273 2732 2337
rect 2748 2333 2812 2337
rect 2828 2333 2892 2337
rect 2748 2277 2786 2333
rect 2786 2277 2812 2333
rect 2828 2277 2842 2333
rect 2842 2277 2892 2333
rect 2748 2273 2812 2277
rect 2828 2273 2892 2277
rect 2908 2273 2972 2337
rect 2988 2333 3052 2337
rect 2988 2277 3010 2333
rect 3010 2277 3052 2333
rect 2988 2273 3052 2277
rect 3068 2273 3132 2337
rect 3148 2273 3212 2337
rect 3228 2333 3292 2337
rect 3228 2277 3234 2333
rect 3234 2277 3290 2333
rect 3290 2277 3292 2333
rect 3228 2273 3292 2277
rect 3308 2273 3372 2337
rect 3388 2273 3452 2337
rect 3468 2333 3532 2337
rect 3468 2277 3514 2333
rect 3514 2277 3532 2333
rect 3468 2273 3532 2277
rect 3548 2273 3612 2337
rect 3628 2333 3692 2337
rect 3708 2333 3772 2337
rect 3628 2277 3682 2333
rect 3682 2277 3692 2333
rect 3708 2277 3738 2333
rect 3738 2277 3772 2333
rect 3628 2273 3692 2277
rect 3708 2273 3772 2277
rect 3788 2273 3852 2337
rect 3868 2333 3932 2337
rect 3948 2333 4012 2337
rect 3868 2277 3906 2333
rect 3906 2277 3932 2333
rect 3948 2277 3962 2333
rect 3962 2277 4012 2333
rect 3868 2273 3932 2277
rect 3948 2273 4012 2277
rect 4028 2273 4092 2337
rect 4108 2333 4172 2337
rect 4108 2277 4130 2333
rect 4130 2277 4172 2333
rect 4108 2273 4172 2277
rect 4188 2273 4252 2337
rect 4268 2273 4332 2337
rect 4348 2273 4412 2337
rect 28 61 92 65
rect 28 5 42 61
rect 42 5 92 61
rect 28 1 92 5
rect 108 1 172 65
rect 188 1 252 65
rect 268 61 332 65
rect 268 5 322 61
rect 322 5 332 61
rect 268 1 332 5
rect 348 1 412 65
rect 428 61 492 65
rect 508 61 572 65
rect 428 5 490 61
rect 490 5 492 61
rect 508 5 546 61
rect 546 5 572 61
rect 428 1 492 5
rect 508 1 572 5
rect 588 1 652 65
rect 668 61 732 65
rect 748 61 812 65
rect 668 5 714 61
rect 714 5 732 61
rect 748 5 770 61
rect 770 5 812 61
rect 668 1 732 5
rect 748 1 812 5
rect 828 1 892 65
rect 908 61 972 65
rect 988 61 1052 65
rect 908 5 938 61
rect 938 5 972 61
rect 988 5 994 61
rect 994 5 1052 61
rect 908 1 972 5
rect 988 1 1052 5
rect 1068 1 1132 65
rect 1148 61 1212 65
rect 1148 5 1162 61
rect 1162 5 1212 61
rect 1148 1 1212 5
rect 1228 1 1292 65
rect 1308 1 1372 65
rect 1388 61 1452 65
rect 1388 5 1442 61
rect 1442 5 1452 61
rect 1388 1 1452 5
rect 1468 1 1532 65
rect 1548 61 1612 65
rect 1628 61 1692 65
rect 1548 5 1610 61
rect 1610 5 1612 61
rect 1628 5 1666 61
rect 1666 5 1692 61
rect 1548 1 1612 5
rect 1628 1 1692 5
rect 1708 1 1772 65
rect 1788 61 1852 65
rect 1868 61 1932 65
rect 1788 5 1834 61
rect 1834 5 1852 61
rect 1868 5 1890 61
rect 1890 5 1932 61
rect 1788 1 1852 5
rect 1868 1 1932 5
rect 1948 1 2012 65
rect 2028 61 2092 65
rect 2108 61 2172 65
rect 2028 5 2058 61
rect 2058 5 2092 61
rect 2108 5 2114 61
rect 2114 5 2172 61
rect 2028 1 2092 5
rect 2108 1 2172 5
rect 2188 1 2252 65
rect 2268 61 2332 65
rect 2268 5 2282 61
rect 2282 5 2332 61
rect 2268 1 2332 5
rect 2348 1 2412 65
rect 2428 1 2492 65
rect 2508 61 2572 65
rect 2508 5 2562 61
rect 2562 5 2572 61
rect 2508 1 2572 5
rect 2588 1 2652 65
rect 2668 61 2732 65
rect 2748 61 2812 65
rect 2668 5 2730 61
rect 2730 5 2732 61
rect 2748 5 2786 61
rect 2786 5 2812 61
rect 2668 1 2732 5
rect 2748 1 2812 5
rect 2828 1 2892 65
rect 2908 61 2972 65
rect 2988 61 3052 65
rect 2908 5 2954 61
rect 2954 5 2972 61
rect 2988 5 3010 61
rect 3010 5 3052 61
rect 2908 1 2972 5
rect 2988 1 3052 5
rect 3068 1 3132 65
rect 3148 61 3212 65
rect 3228 61 3292 65
rect 3148 5 3178 61
rect 3178 5 3212 61
rect 3228 5 3234 61
rect 3234 5 3292 61
rect 3148 1 3212 5
rect 3228 1 3292 5
rect 3308 1 3372 65
rect 3388 61 3452 65
rect 3388 5 3402 61
rect 3402 5 3452 61
rect 3388 1 3452 5
rect 3468 1 3532 65
rect 3548 1 3612 65
rect 3628 61 3692 65
rect 3628 5 3682 61
rect 3682 5 3692 61
rect 3628 1 3692 5
rect 3708 1 3772 65
rect 3788 61 3852 65
rect 3868 61 3932 65
rect 3788 5 3850 61
rect 3850 5 3852 61
rect 3868 5 3906 61
rect 3906 5 3932 61
rect 3788 1 3852 5
rect 3868 1 3932 5
rect 3948 1 4012 65
rect 4028 61 4092 65
rect 4108 61 4172 65
rect 4028 5 4074 61
rect 4074 5 4092 61
rect 4108 5 4130 61
rect 4130 5 4172 61
rect 4028 1 4092 5
rect 4108 1 4172 5
rect 4188 1 4252 65
rect 4268 61 4332 65
rect 4348 61 4412 65
rect 4268 5 4298 61
rect 4298 5 4332 61
rect 4348 5 4354 61
rect 4354 5 4412 61
rect 4268 1 4332 5
rect 4348 1 4412 5
<< metal4 >>
rect 0 2337 4498 2338
rect 0 2273 28 2337
rect 92 2273 108 2337
rect 172 2273 188 2337
rect 252 2273 268 2337
rect 332 2273 348 2337
rect 412 2273 428 2337
rect 492 2273 508 2337
rect 572 2273 588 2337
rect 652 2273 668 2337
rect 732 2273 748 2337
rect 812 2273 828 2337
rect 892 2273 908 2337
rect 972 2273 988 2337
rect 1052 2273 1068 2337
rect 1132 2273 1148 2337
rect 1212 2273 1228 2337
rect 1292 2273 1308 2337
rect 1372 2273 1388 2337
rect 1452 2273 1468 2337
rect 1532 2273 1548 2337
rect 1612 2273 1628 2337
rect 1692 2273 1708 2337
rect 1772 2273 1788 2337
rect 1852 2273 1868 2337
rect 1932 2273 1948 2337
rect 2012 2273 2028 2337
rect 2092 2273 2108 2337
rect 2172 2273 2188 2337
rect 2252 2273 2268 2337
rect 2332 2273 2348 2337
rect 2412 2273 2428 2337
rect 2492 2273 2508 2337
rect 2572 2273 2588 2337
rect 2652 2273 2668 2337
rect 2732 2273 2748 2337
rect 2812 2273 2828 2337
rect 2892 2273 2908 2337
rect 2972 2273 2988 2337
rect 3052 2273 3068 2337
rect 3132 2273 3148 2337
rect 3212 2273 3228 2337
rect 3292 2273 3308 2337
rect 3372 2273 3388 2337
rect 3452 2273 3468 2337
rect 3532 2273 3548 2337
rect 3612 2273 3628 2337
rect 3692 2273 3708 2337
rect 3772 2273 3788 2337
rect 3852 2273 3868 2337
rect 3932 2273 3948 2337
rect 4012 2273 4028 2337
rect 4092 2273 4108 2337
rect 4172 2273 4188 2337
rect 4252 2273 4268 2337
rect 4332 2273 4348 2337
rect 4412 2273 4498 2337
rect 0 2272 4498 2273
rect 120 2263 420 2272
rect 0 66 60 2212
rect 120 2027 152 2263
rect 388 2027 420 2263
rect 120 126 180 2027
rect 240 311 300 1967
rect 360 371 420 2027
rect 480 311 540 2212
rect 240 75 272 311
rect 508 75 540 311
rect 600 126 660 2272
rect 240 66 540 75
rect 720 66 780 2212
rect 840 126 900 2272
rect 960 66 1020 2212
rect 1080 126 1140 2272
rect 1200 66 1260 2212
rect 1320 126 1380 2272
rect 1560 2263 1860 2272
rect 1440 66 1500 2212
rect 1560 2027 1592 2263
rect 1828 2027 1860 2263
rect 1560 126 1620 2027
rect 1680 311 1740 1967
rect 1800 371 1860 2027
rect 1920 311 1980 2212
rect 1680 75 1712 311
rect 1948 75 1980 311
rect 2040 126 2100 2272
rect 1680 66 1980 75
rect 2160 66 2220 2212
rect 2280 126 2340 2272
rect 2400 66 2460 2212
rect 2520 126 2580 2272
rect 2640 66 2700 2212
rect 2760 126 2820 2272
rect 3000 2263 3300 2272
rect 2880 66 2940 2212
rect 3000 2027 3032 2263
rect 3268 2027 3300 2263
rect 3000 126 3060 2027
rect 3120 311 3180 1967
rect 3240 371 3300 2027
rect 3360 311 3420 2212
rect 3120 75 3152 311
rect 3388 75 3420 311
rect 3480 126 3540 2272
rect 3120 66 3420 75
rect 3600 66 3660 2212
rect 3720 126 3780 2272
rect 3840 66 3900 2212
rect 3960 126 4020 2272
rect 4080 66 4140 2212
rect 4200 126 4260 2272
rect 4320 66 4498 2212
rect 0 65 4498 66
rect 0 1 28 65
rect 92 1 108 65
rect 172 1 188 65
rect 252 1 268 65
rect 332 1 348 65
rect 412 1 428 65
rect 492 1 508 65
rect 572 1 588 65
rect 652 1 668 65
rect 732 1 748 65
rect 812 1 828 65
rect 892 1 908 65
rect 972 1 988 65
rect 1052 1 1068 65
rect 1132 1 1148 65
rect 1212 1 1228 65
rect 1292 1 1308 65
rect 1372 1 1388 65
rect 1452 1 1468 65
rect 1532 1 1548 65
rect 1612 1 1628 65
rect 1692 1 1708 65
rect 1772 1 1788 65
rect 1852 1 1868 65
rect 1932 1 1948 65
rect 2012 1 2028 65
rect 2092 1 2108 65
rect 2172 1 2188 65
rect 2252 1 2268 65
rect 2332 1 2348 65
rect 2412 1 2428 65
rect 2492 1 2508 65
rect 2572 1 2588 65
rect 2652 1 2668 65
rect 2732 1 2748 65
rect 2812 1 2828 65
rect 2892 1 2908 65
rect 2972 1 2988 65
rect 3052 1 3068 65
rect 3132 1 3148 65
rect 3212 1 3228 65
rect 3292 1 3308 65
rect 3372 1 3388 65
rect 3452 1 3468 65
rect 3532 1 3548 65
rect 3612 1 3628 65
rect 3692 1 3708 65
rect 3772 1 3788 65
rect 3852 1 3868 65
rect 3932 1 3948 65
rect 4012 1 4028 65
rect 4092 1 4108 65
rect 4172 1 4188 65
rect 4252 1 4268 65
rect 4332 1 4348 65
rect 4412 1 4498 65
rect 0 0 4498 1
<< via4 >>
rect 152 2027 388 2263
rect 272 75 508 311
rect 1592 2027 1828 2263
rect 1712 75 1948 311
rect 3032 2027 3268 2263
rect 3152 75 3388 311
<< metal5 >>
rect 0 2263 4498 2338
rect 0 2027 152 2263
rect 388 2027 1592 2263
rect 1828 2027 3032 2263
rect 3268 2027 4498 2263
rect 0 2003 4498 2027
rect 0 655 320 2003
rect 640 335 960 1683
rect 1280 655 1600 2003
rect 1920 335 2240 1683
rect 2560 655 2880 2003
rect 3200 335 3520 1683
rect 3840 655 4498 2003
rect 0 311 4498 335
rect 0 75 272 311
rect 508 75 1712 311
rect 1948 75 3152 311
rect 3388 75 4498 311
rect 0 0 4498 75
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 1294370
string GDS_START 1231582
<< end >>
