magic
tech sky130A
timestamp 1634425727
<< pwell >>
rect -148 -465 148 465
<< nmoslvt >>
rect -50 260 50 360
rect -50 105 50 205
rect -50 -50 50 50
rect -50 -205 50 -105
rect -50 -360 50 -260
<< ndiff >>
rect -79 354 -50 360
rect -79 266 -73 354
rect -56 266 -50 354
rect -79 260 -50 266
rect 50 354 79 360
rect 50 266 56 354
rect 73 266 79 354
rect 50 260 79 266
rect -79 199 -50 205
rect -79 111 -73 199
rect -56 111 -50 199
rect -79 105 -50 111
rect 50 199 79 205
rect 50 111 56 199
rect 73 111 79 199
rect 50 105 79 111
rect -79 44 -50 50
rect -79 -44 -73 44
rect -56 -44 -50 44
rect -79 -50 -50 -44
rect 50 44 79 50
rect 50 -44 56 44
rect 73 -44 79 44
rect 50 -50 79 -44
rect -79 -111 -50 -105
rect -79 -199 -73 -111
rect -56 -199 -50 -111
rect -79 -205 -50 -199
rect 50 -111 79 -105
rect 50 -199 56 -111
rect 73 -199 79 -111
rect 50 -205 79 -199
rect -79 -266 -50 -260
rect -79 -354 -73 -266
rect -56 -354 -50 -266
rect -79 -360 -50 -354
rect 50 -266 79 -260
rect 50 -354 56 -266
rect 73 -354 79 -266
rect 50 -360 79 -354
<< ndiffc >>
rect -73 266 -56 354
rect 56 266 73 354
rect -73 111 -56 199
rect 56 111 73 199
rect -73 -44 -56 44
rect 56 -44 73 44
rect -73 -199 -56 -111
rect 56 -199 73 -111
rect -73 -354 -56 -266
rect 56 -354 73 -266
<< psubdiff >>
rect -130 430 -82 447
rect 82 430 130 447
rect -130 399 -113 430
rect 113 399 130 430
<< psubdiffcont >>
rect -82 430 82 447
<< poly >>
rect -50 396 50 404
rect -50 379 -42 396
rect 42 379 50 396
rect -50 360 50 379
rect -50 241 50 260
rect -50 224 -42 241
rect 42 224 50 241
rect -50 205 50 224
rect -50 86 50 105
rect -50 69 -42 86
rect 42 69 50 86
rect -50 50 50 69
rect -50 -69 50 -50
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -50 -105 50 -86
rect -50 -224 50 -205
rect -50 -241 -42 -224
rect 42 -241 50 -224
rect -50 -260 50 -241
rect -50 -379 50 -360
rect -50 -396 -42 -379
rect 42 -396 50 -379
rect -50 -404 50 -396
<< polycont >>
rect -42 379 42 396
rect -42 224 42 241
rect -42 69 42 86
rect -42 -86 42 -69
rect -42 -241 42 -224
rect -42 -396 42 -379
<< locali >>
rect -130 430 -82 447
rect 82 430 130 447
rect -130 399 -113 430
rect 113 399 130 430
rect -50 379 -42 396
rect 42 379 50 396
rect -73 354 -56 362
rect -73 258 -56 266
rect 56 354 73 362
rect 56 258 73 266
rect -50 224 -42 241
rect 42 224 50 241
rect -73 199 -56 207
rect -73 103 -56 111
rect 56 199 73 207
rect 56 103 73 111
rect -50 69 -42 86
rect 42 69 50 86
rect -73 44 -56 52
rect -73 -52 -56 -44
rect 56 44 73 52
rect 56 -52 73 -44
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -73 -111 -56 -103
rect -73 -207 -56 -199
rect 56 -111 73 -103
rect 56 -207 73 -199
rect -50 -241 -42 -224
rect 42 -241 50 -224
rect -73 -266 -56 -258
rect -73 -362 -56 -354
rect 56 -266 73 -258
rect 56 -362 73 -354
rect -50 -396 -42 -379
rect 42 -396 50 -379
<< viali >>
rect -42 379 42 396
rect -73 266 -56 354
rect 56 266 73 354
rect -42 224 42 241
rect -73 111 -56 199
rect 56 111 73 199
rect -42 69 42 86
rect -73 -44 -56 44
rect 56 -44 73 44
rect -42 -86 42 -69
rect -73 -199 -56 -111
rect 56 -199 73 -111
rect -42 -241 42 -224
rect -73 -354 -56 -266
rect 56 -354 73 -266
rect -42 -396 42 -379
<< metal1 >>
rect 7 399 78 400
rect -48 396 78 399
rect -48 379 -42 396
rect 42 379 78 396
rect -48 376 78 379
rect 7 375 78 376
rect -76 354 -53 360
rect -76 266 -73 354
rect -56 266 -53 354
rect 52 354 77 375
rect 52 329 56 354
rect -76 260 -53 266
rect 53 266 56 329
rect 73 329 77 354
rect 73 266 76 329
rect 53 260 76 266
rect 39 245 75 246
rect 39 244 76 245
rect -48 241 76 244
rect -48 224 -42 241
rect 42 224 76 241
rect -48 221 76 224
rect -76 199 -53 205
rect 51 199 76 221
rect -76 111 -73 199
rect -56 111 -53 199
rect -76 105 -53 111
rect 53 111 56 199
rect 73 111 76 199
rect 53 105 76 111
rect -48 86 49 89
rect -48 69 -42 86
rect 42 69 49 86
rect -48 66 49 69
rect -76 44 -53 50
rect -76 -44 -73 44
rect -56 -44 -53 44
rect -76 -50 -53 -44
rect 53 44 76 50
rect 53 -44 56 44
rect 73 -44 76 44
rect 53 -50 76 -44
rect -48 -68 48 -66
rect -48 -69 76 -68
rect -48 -86 -42 -69
rect 42 -86 76 -69
rect -48 -89 76 -86
rect -76 -111 -53 -105
rect -76 -199 -73 -111
rect -56 -199 -53 -111
rect 51 -111 76 -89
rect 51 -114 56 -111
rect -76 -205 -53 -199
rect 53 -199 56 -114
rect 73 -199 76 -111
rect 53 -205 76 -199
rect -48 -222 48 -221
rect -48 -224 76 -222
rect -48 -241 -42 -224
rect 42 -241 76 -224
rect -48 -244 76 -241
rect -76 -266 -53 -260
rect -76 -354 -73 -266
rect -56 -354 -53 -266
rect 52 -266 76 -244
rect 52 -271 56 -266
rect -76 -360 -53 -354
rect 53 -354 56 -271
rect 73 -354 76 -266
rect 53 -360 76 -354
rect -48 -379 48 -376
rect -48 -396 -42 -379
rect 42 -396 48 -379
rect -48 -399 48 -396
<< labels >>
flabel nmoslvt -50 -50 50 50 0 FreeSans 240 0 0 0 M18,17
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -121 -438 121 438
string parameters w 1 l 1 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
