magic
tech sky130A
timestamp 1634658360
<< metal1 >>
rect -697 773 -640 781
rect -395 779 -280 816
rect 257 797 390 811
rect -536 773 -280 779
rect -697 75 -652 773
rect -536 700 -391 773
rect -316 700 -280 773
rect -536 681 -280 700
rect -395 670 -280 681
rect -402 625 -287 650
rect -532 622 -287 625
rect -532 555 -391 622
rect -535 549 -391 555
rect -316 549 -287 622
rect -535 527 -287 549
rect -535 511 -503 527
rect -565 485 -503 511
rect -402 504 -287 527
rect -537 463 -94 470
rect -537 389 -192 463
rect -108 389 -94 463
rect -537 372 -94 389
rect -389 314 -290 317
rect -533 301 -290 314
rect -533 228 -391 301
rect -316 228 -290 301
rect -533 216 -290 228
rect -389 215 -290 216
rect -398 160 -283 183
rect -698 -293 -652 75
rect -536 151 -283 160
rect -536 78 -392 151
rect -317 78 -283 151
rect -536 62 -283 78
rect -398 37 -283 62
rect -698 -834 -654 -293
rect -15 -639 30 790
rect 257 781 289 797
rect 146 700 289 781
rect 377 781 390 797
rect 377 700 395 781
rect 146 681 395 700
rect 257 677 390 681
rect 257 640 390 659
rect 257 625 287 640
rect 146 568 287 625
rect 143 543 287 568
rect 375 625 390 640
rect 375 543 395 625
rect 143 526 395 543
rect 149 510 174 526
rect 188 525 395 526
rect 138 486 174 510
rect 146 460 534 470
rect 146 389 440 460
rect 524 389 534 460
rect 146 370 534 389
rect 259 369 534 370
rect 261 324 394 347
rect 261 315 282 324
rect 145 227 282 315
rect 370 227 394 324
rect 145 215 394 227
rect 261 214 394 215
rect 148 162 149 175
rect 266 165 394 178
rect 266 162 279 165
rect 148 96 279 162
rect 143 68 279 96
rect 367 68 394 165
rect 143 62 394 68
rect 143 58 178 62
rect 133 22 178 58
rect 266 38 394 62
rect 143 20 178 22
rect 648 -376 683 797
rect 932 784 1037 795
rect 932 775 954 784
rect 798 700 954 775
rect 1023 700 1037 784
rect 798 681 1037 700
rect 798 677 937 681
rect 796 612 1039 621
rect 796 530 944 612
rect 804 505 827 530
rect 844 529 944 530
rect 1021 529 1039 612
rect 844 523 1039 529
rect 795 483 827 505
rect 927 466 1201 469
rect 799 461 1201 466
rect 799 374 1119 461
rect 1182 374 1201 461
rect 799 365 1201 374
rect 803 301 1046 311
rect 803 218 950 301
rect 1027 218 1046 301
rect 803 213 1046 218
rect 802 153 1045 156
rect 802 107 947 153
rect 799 70 947 107
rect 1024 70 1045 153
rect 799 58 1045 70
rect 799 50 832 58
rect 783 18 832 50
rect 783 14 828 18
rect 1286 -186 1329 805
rect 1447 774 1714 780
rect 1447 688 1619 774
rect 1699 688 1714 774
rect 1447 680 1714 688
rect 1440 621 1707 625
rect 1440 571 1610 621
rect 1439 535 1610 571
rect 1690 535 1707 621
rect 1439 526 1707 535
rect 1447 508 1472 526
rect 1492 525 1707 526
rect 1444 485 1474 508
rect 1444 458 1976 471
rect 1444 383 1866 458
rect 1950 383 1976 458
rect 1444 368 1976 383
rect 1444 312 1711 315
rect 1444 226 1623 312
rect 1703 226 1711 312
rect 1444 215 1711 226
rect 1416 176 1442 196
rect 1442 151 1709 158
rect 1442 111 1610 151
rect 1441 65 1610 111
rect 1690 65 1709 151
rect 1441 59 1709 65
rect 1448 43 1471 59
rect 1488 58 1709 59
rect 1425 26 1434 42
rect 1443 20 1475 43
rect 1286 -196 1504 -186
rect 1286 -205 2210 -196
rect 1286 -306 2100 -205
rect 2189 -306 2210 -205
rect 1286 -321 2210 -306
rect 1315 -323 2210 -321
rect 648 -380 822 -376
rect 648 -412 1981 -380
rect 648 -534 1860 -412
rect 1955 -534 1981 -412
rect 648 -552 1981 -534
rect 648 -555 822 -552
rect -15 -640 151 -639
rect -15 -661 1214 -640
rect -15 -756 1101 -661
rect 1202 -756 1214 -661
rect -15 -769 1214 -756
rect 196 -780 1214 -769
rect -630 -834 550 -833
rect -698 -851 550 -834
rect -698 -975 461 -851
rect 544 -975 550 -851
rect -698 -996 550 -975
rect -698 -999 -343 -996
<< via1 >>
rect -391 700 -316 773
rect -391 549 -316 622
rect -192 389 -108 463
rect -391 228 -316 301
rect -392 78 -317 151
rect 289 700 377 797
rect 287 543 375 640
rect 440 389 524 460
rect 282 227 370 324
rect 279 68 367 165
rect 954 700 1023 784
rect 944 529 1021 612
rect 1119 374 1182 461
rect 950 218 1027 301
rect 947 70 1024 153
rect 1619 688 1699 774
rect 1610 535 1690 621
rect 1866 383 1950 458
rect 1623 226 1703 312
rect 1610 65 1690 151
rect 2100 -306 2189 -205
rect 1860 -534 1955 -412
rect 1101 -756 1202 -661
rect 461 -975 544 -851
<< metal2 >>
rect -426 926 -246 1429
rect -205 932 -71 1022
rect -402 773 -264 926
rect -402 700 -391 773
rect -316 700 -264 773
rect -402 622 -264 700
rect -402 549 -391 622
rect -316 549 -264 622
rect -402 301 -264 549
rect -402 228 -391 301
rect -316 228 -264 301
rect -402 151 -264 228
rect -402 78 -392 151
rect -317 78 -264 151
rect -402 -107 -264 78
rect -204 463 -66 932
rect 251 829 399 1414
rect -204 389 -192 463
rect -108 389 -66 463
rect -204 -107 -66 389
rect 259 797 397 829
rect 259 700 289 797
rect 377 700 397 797
rect 259 640 397 700
rect 259 543 287 640
rect 375 543 397 640
rect 259 324 397 543
rect 435 460 554 932
rect 925 867 1049 1420
rect 1596 932 1747 1408
rect 2067 1055 2248 1532
rect 435 389 440 460
rect 524 389 554 460
rect 927 784 1046 867
rect 927 700 954 784
rect 1023 700 1046 784
rect 927 612 1046 700
rect 927 529 944 612
rect 1021 529 1046 612
rect 259 227 282 324
rect 370 227 397 324
rect 259 165 397 227
rect 259 68 279 165
rect 367 68 397 165
rect 259 -107 397 68
rect -204 -409 -70 -107
rect 436 -134 553 389
rect 927 301 1046 529
rect 927 218 950 301
rect 1027 218 1046 301
rect 927 153 1046 218
rect 927 70 947 153
rect 1024 70 1046 153
rect 927 -107 1046 70
rect 1099 461 1218 932
rect 1099 374 1119 461
rect 1182 374 1218 461
rect 1099 -94 1218 374
rect 1091 -134 1218 -94
rect 1595 774 1759 932
rect 1595 688 1619 774
rect 1699 688 1759 774
rect 1595 621 1759 688
rect 1595 535 1610 621
rect 1690 535 1759 621
rect 1595 312 1759 535
rect 1595 226 1623 312
rect 1703 226 1759 312
rect 1595 151 1759 226
rect 1845 458 2009 932
rect 1845 383 1866 458
rect 1950 383 2009 458
rect 1845 154 2009 383
rect 1595 65 1610 151
rect 1690 65 1759 151
rect 1595 -107 1759 65
rect 1842 152 2009 154
rect 1842 -94 1999 152
rect -215 -1345 -64 -409
rect 437 -851 550 -134
rect 1095 -661 1211 -134
rect 1839 -151 1999 -94
rect 1842 -412 1999 -151
rect 1842 -534 1860 -412
rect 1955 -534 1999 -412
rect 2076 -205 2248 1055
rect 2076 -306 2100 -205
rect 2189 -306 2248 -205
rect 2076 -492 2248 -306
rect 1842 -552 1999 -534
rect 1095 -756 1101 -661
rect 1202 -756 1211 -661
rect 1095 -815 1211 -756
rect 437 -975 461 -851
rect 544 -975 550 -851
rect 437 -990 550 -975
rect -641 -1494 -61 -1345
use sky130_fd_pr__nfet_01v8_lvt_M15_14  M15_14
timestamp 1634425567
transform 1 0 751 0 1 416
box -148 -465 148 465
use sky130_fd_pr__nfet_01v8_lvt_M18_17  M18_17
timestamp 1634425727
transform 1 0 1395 0 1 419
box -148 -465 148 465
use sky130_fd_pr__nfet_01v8_lvt_M6_7  M6_7
timestamp 1634425503
transform 1 0 97 0 1 420
box -148 -465 148 465
use sky130_fd_pr__nfet_01v8_lvt_M4_5  M4_5
timestamp 1634457025
transform 1 0 -582 0 1 420
box -148 -465 148 465
<< labels >>
flabel metal2 2076 -205 2248 1173 0 FreeSans 400 0 0 0 DM18
flabel space -1344 -1494 -61 -1345 0 FreeSans 400 0 0 0 SM4
flabel metal1 1315 -323 2100 -196 0 FreeSans 400 0 0 0 DM18
flabel metal1 648 -552 1860 -380 0 FreeSans 400 0 0 0 DM15
flabel metal1 196 -780 1101 -640 0 FreeSans 400 0 0 0 DM6
flabel metal1 -15 -769 30 790 0 FreeSans 400 0 0 0 DM6
flabel metal1 648 -555 683 797 0 FreeSans 400 0 0 0 DM15
flabel metal1 1286 -321 1329 805 0 FreeSans 400 0 0 0 DM18
flabel metal2 1595 312 1759 535 0 FreeSans 400 0 0 0 DM17
flabel metal2 -316 -107 -264 1429 0 FreeSans 400 0 0 0 DM5
flabel metal2 -402 622 -264 700 0 FreeSans 400 0 0 0 DM5
flabel metal2 251 829 399 1414 0 FreeSans 400 0 0 0 DM7
flabel via1 287 543 375 640 0 FreeSans 400 0 0 0 DM7
flabel metal1 -630 -996 461 -833 0 FreeSans 400 0 0 0 SM6
flabel metal1 -697 -293 -652 781 0 FreeSans 400 0 0 0 SM6
flabel metal1 -697 -293 -690 -291 0 FreeSans 400 0 0 0 SM6
flabel metal2 1099 -134 1218 374 0 FreeSans 400 0 0 0 SM15
flabel metal2 927 612 1046 700 0 FreeSans 400 0 0 0 DM14
<< end >>
