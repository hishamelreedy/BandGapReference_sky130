magic
tech sky130A
timestamp 1634058968
<< nwell >>
rect -97 -81 97 81
<< pmoslvt >>
rect -50 -50 50 50
<< pdiff >>
rect -79 44 -50 50
rect -79 -44 -73 44
rect -56 -44 -50 44
rect -79 -50 -50 -44
rect 50 44 79 50
rect 50 -44 56 44
rect 73 -44 79 44
rect 50 -50 79 -44
<< pdiffc >>
rect -73 -44 -56 44
rect 56 -44 73 44
<< poly >>
rect -50 50 50 63
rect -50 -63 50 -50
<< locali >>
rect -73 44 -56 52
rect -73 -52 -56 -44
rect 56 44 73 52
rect 56 -52 73 -44
<< viali >>
rect -73 -44 -56 44
rect 56 -44 73 44
<< metal1 >>
rect -76 44 -53 50
rect -76 -44 -73 44
rect -56 -44 -53 44
rect -76 -50 -53 -44
rect 53 44 76 50
rect 53 -44 56 44
rect 73 -44 76 44
rect 53 -50 76 -44
<< labels >>
flabel nwell -97 -81 97 81 0 FreeSans 400 0 0 0 M11
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 1 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
