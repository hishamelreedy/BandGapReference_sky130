magic
tech sky130A
magscale 1 2
timestamp 1634658069
<< metal1 >>
rect -2156 5126 -2012 5138
rect -2156 5034 -2142 5126
rect -2028 5034 -2012 5126
rect -2156 5020 -2012 5034
rect -1412 5130 -1264 5160
rect -1412 5042 -1390 5130
rect -1294 5042 -1264 5130
rect -1412 5026 -1264 5042
rect -884 5146 -732 5174
rect -884 5054 -868 5146
rect -766 5054 -732 5146
rect -1392 5024 -1276 5026
rect -884 5024 -732 5054
rect -382 5150 -228 5168
rect -382 5058 -362 5150
rect -258 5058 -228 5150
rect -382 5038 -228 5058
rect 320 5136 512 5150
rect 320 5038 346 5136
rect 498 5038 512 5136
rect -2392 4716 -2294 4728
rect -2392 4646 -2382 4716
rect -2304 4646 -2294 4716
rect -2392 4630 -2294 4646
rect -3014 4230 -2930 4238
rect -3014 4170 -3004 4230
rect -2942 4170 -2930 4230
rect -3014 4014 -2930 4170
rect -2996 3596 -2958 4014
rect -2360 3608 -2324 4630
rect -2106 3570 -2058 5020
rect -1878 4714 -1758 4728
rect -1878 4638 -1852 4714
rect -1782 4638 -1758 4714
rect -1878 4616 -1758 4638
rect -1842 3568 -1806 4616
rect -1360 3574 -1308 5024
rect -1182 4196 -952 4234
rect -1182 4098 -1154 4196
rect -1044 4098 -952 4196
rect -1182 4012 -952 4098
rect -1106 3008 -1038 4012
rect -844 3594 -788 5024
rect -700 4204 -432 4248
rect -700 4088 -592 4204
rect -448 4088 -432 4204
rect -700 4076 -432 4088
rect -698 3998 -432 4076
rect -598 3030 -530 3998
rect -330 3584 -276 5038
rect 320 5024 512 5038
rect 80 4748 244 4772
rect 80 4642 106 4748
rect 226 4642 244 4748
rect 80 4630 244 4642
rect 126 3582 184 4630
rect 392 3578 440 5024
rect 590 4708 760 4720
rect 590 4618 618 4708
rect 740 4618 760 4708
rect 590 4614 760 4618
rect 646 3566 704 4614
rect 968 4030 1446 4032
rect 968 4024 1448 4030
rect 968 3934 994 4024
rect 1094 3934 1448 4024
rect 968 3922 1448 3934
rect 1410 3600 1448 3922
rect -3268 2008 -3208 2130
rect -2730 2120 -2710 2126
rect -3272 1982 -3154 2008
rect -3272 1914 -3028 1982
rect -3196 1218 -3028 1914
rect -2934 1978 -2766 1980
rect -2734 1978 -2704 2120
rect 1158 2060 1180 2108
rect 1158 2044 1186 2060
rect -2934 1950 -2704 1978
rect -2934 1934 -2706 1950
rect -2934 1236 -2766 1934
rect -2298 1600 -2118 1986
rect -2034 1742 -1874 1982
rect -1274 1600 -1122 1992
rect -1024 1600 -872 1992
rect -764 1600 -612 1994
rect 1158 1990 1194 2044
rect 1674 2028 1700 2080
rect -508 1600 -352 1966
rect 200 1600 378 1982
rect 458 1600 636 1982
rect 1158 1946 1378 1990
rect 1162 1942 1378 1946
rect -2298 1574 660 1600
rect -2288 1374 660 1574
rect 1212 1380 1378 1942
rect -3216 1016 -3006 1218
rect -3216 886 -3202 1016
rect -3026 886 -3006 1016
rect -2946 1016 -2748 1236
rect 1202 1084 1378 1380
rect 1212 1024 1378 1084
rect -2946 926 -2922 1016
rect -2784 926 -2748 1016
rect -2946 924 -2748 926
rect 1206 1008 1384 1024
rect -3216 822 -3006 886
rect 1206 882 1232 1008
rect 1366 882 1384 1008
rect 1206 832 1384 882
rect 1482 974 1616 2012
rect 1674 1990 1704 2028
rect 1626 1966 1704 1990
rect 1626 1962 1702 1966
rect 1482 834 1506 974
rect 1596 834 1616 974
rect 1482 830 1616 834
<< via1 >>
rect -2142 5034 -2028 5126
rect -1390 5042 -1294 5130
rect -868 5054 -766 5146
rect -362 5058 -258 5150
rect 346 5038 498 5136
rect -2382 4646 -2304 4716
rect -3004 4170 -2942 4230
rect -1852 4638 -1782 4714
rect -1154 4098 -1044 4196
rect -592 4088 -448 4204
rect 106 4642 226 4748
rect 618 4618 740 4708
rect 994 3934 1094 4024
rect -3202 886 -3026 1016
rect -2922 926 -2784 1016
rect 1232 882 1366 1008
rect 1506 834 1596 974
<< metal2 >>
rect -3406 5150 1200 5224
rect -3406 5146 -362 5150
rect -3406 5130 -868 5146
rect -3406 5126 -1390 5130
rect -3406 5034 -2142 5126
rect -2028 5042 -1390 5126
rect -1294 5054 -868 5130
rect -766 5058 -362 5146
rect -258 5136 1200 5150
rect -258 5058 346 5136
rect -766 5054 346 5058
rect -1294 5042 346 5054
rect -2028 5038 346 5042
rect 498 5038 1200 5136
rect -2028 5034 1200 5038
rect -3406 5010 1200 5034
rect -3410 4748 1200 4820
rect -3410 4716 106 4748
rect -3410 4646 -2382 4716
rect -2304 4714 106 4716
rect -2304 4646 -1852 4714
rect -3410 4638 -1852 4646
rect -1782 4642 106 4714
rect 226 4708 1200 4748
rect 226 4642 618 4708
rect -1782 4638 618 4642
rect -3410 4618 618 4638
rect 740 4618 1200 4708
rect -3410 4606 1200 4618
rect -2662 4278 -2398 4290
rect -3458 4230 -1760 4278
rect -3458 4170 -3004 4230
rect -2942 4170 -1760 4230
rect -3458 4152 -1760 4170
rect -1686 4228 -1430 4284
rect -244 4236 6 4276
rect -2662 3958 -2398 4152
rect -1686 4092 -1638 4228
rect -1474 4204 -1430 4228
rect -338 4234 32 4236
rect -602 4208 -434 4212
rect -338 4208 -192 4234
rect -602 4204 -192 4208
rect -1474 4196 -1030 4204
rect -1474 4098 -1154 4196
rect -1044 4098 -1030 4196
rect -1474 4092 -1030 4098
rect -1686 4000 -1430 4092
rect -602 4088 -592 4204
rect -448 4088 -192 4204
rect -602 4076 -192 4088
rect -338 4072 -192 4076
rect -30 4072 32 4234
rect -338 4064 32 4072
rect -244 4038 6 4064
rect 824 4042 944 4062
rect 824 4024 1116 4042
rect -2662 3946 -2372 3958
rect 824 3946 994 4024
rect -2662 3934 994 3946
rect 1094 3934 1116 4024
rect -2662 3906 1116 3934
rect -2662 3834 944 3906
rect -2422 3826 944 3834
rect -2422 3812 864 3826
rect -3198 1024 -2980 1030
rect -3490 1016 1910 1024
rect -3490 886 -3202 1016
rect -3026 926 -2922 1016
rect -2784 1014 1910 1016
rect -2784 926 -1650 1014
rect -3026 886 -1650 926
rect -3490 878 -1650 886
rect -1486 1010 1910 1014
rect -1486 880 -208 1010
rect -10 1008 1910 1010
rect -10 882 1232 1008
rect 1366 974 1910 1008
rect 1366 882 1506 974
rect -10 880 1506 882
rect -1486 878 1506 880
rect -3490 834 1506 878
rect 1596 834 1910 974
rect -3490 812 1910 834
rect -3490 810 -3198 812
rect -3024 810 1910 812
<< via2 >>
rect -1638 4092 -1474 4228
rect -192 4072 -30 4234
rect -1650 878 -1486 1014
rect -208 880 -10 1010
<< metal3 >>
rect -222 4268 -8 4270
rect -1672 4228 -1448 4260
rect -1672 4180 -1638 4228
rect -1678 4092 -1638 4180
rect -1474 4092 -1448 4228
rect -1678 4028 -1448 4092
rect -222 4234 -6 4268
rect -222 4072 -192 4234
rect -30 4072 -6 4234
rect -222 4042 -6 4072
rect -1678 1412 -1460 4028
rect -216 1772 -6 4042
rect -1680 1150 -1444 1412
rect -216 1396 -2 1772
rect -1678 1014 -1460 1150
rect -1678 878 -1650 1014
rect -1486 878 -1460 1014
rect -1678 866 -1460 878
rect -216 1100 0 1396
rect -216 1010 -2 1100
rect -216 880 -208 1010
rect -10 880 -2 1010
rect -216 860 -2 880
use sky130_fd_pr__nfet_01v8_lvt_M3  M3_1
timestamp 1634657911
transform 1 0 417 0 1 2816
box -425 -1406 425 1010
use sky130_fd_pr__nfet_01v8_lvt_M3  M3_0
timestamp 1634657911
transform 1 0 -2081 0 1 2818
box -425 -1406 425 1010
use sky130_fd_pr__nfet_01v8_lvt_M2  M2_0
timestamp 1634436918
transform 1 0 -1073 0 1 2830
box -425 -1010 425 1010
use sky130_fd_pr__nfet_01v8_lvt_M1  M1_1
timestamp 1634435886
transform 1 0 -2977 0 1 2808
box -425 -1010 425 1010
use sky130_fd_pr__nfet_01v8_lvt_M1  M1_0
timestamp 1634435886
transform 1 0 1429 0 1 2822
box -425 -1010 425 1010
use sky130_fd_pr__nfet_01v8_lvt_M2  M2_1
timestamp 1634436918
transform 1 0 -557 0 1 2830
box -425 -1010 425 1010
<< labels >>
flabel space -3490 810 2328 1024 0 FreeSans 1600 0 0 0 M1D
flabel metal2 -2942 4152 -1760 4278 0 FreeSans 800 0 0 0 GND
flabel metal2 -10 810 1232 1024 0 FreeSans 1600 0 0 0 M1D
flabel metal2 -1486 810 -208 1024 0 FreeSans 1600 0 0 0 M1D
flabel metal2 -2784 810 -1650 1024 0 FreeSans 1600 0 0 0 M1D
flabel metal2 -3490 810 -3202 1024 0 FreeSans 1600 0 0 0 M1D
flabel space 1596 810 2328 1024 0 FreeSans 1600 0 0 0 M1D
flabel space -3410 4606 2408 4820 0 FreeSans 1600 0 0 0 M3D
flabel space -3406 5010 2412 5224 0 FreeSans 1600 0 0 0 M2D
<< end >>
